
module combined_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7;
  wire   [8:0] carry;

  FADDX1 U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1 U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1 U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR3X1 U1 ( .IN1(A[7]), .IN2(B[7]), .IN3(carry[7]), .Q(DIFF[7]) );
  INVX0 U2 ( .INP(B[1]), .ZN(n7) );
  NAND2X1 U3 ( .IN1(n1), .IN2(B[0]), .QN(carry[1]) );
  INVX0 U4 ( .INP(A[0]), .ZN(n1) );
  INVX0 U5 ( .INP(B[2]), .ZN(n6) );
  INVX0 U6 ( .INP(B[3]), .ZN(n5) );
  INVX0 U7 ( .INP(B[4]), .ZN(n4) );
  INVX0 U8 ( .INP(B[5]), .ZN(n3) );
  INVX0 U9 ( .INP(B[6]), .ZN(n2) );
  XOR2X1 U10 ( .IN1(B[0]), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module combined_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FADDX1 U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XOR3X1 U2_7 ( .IN1(A[7]), .IN2(n2), .IN3(carry[7]), .Q(DIFF[7]) );
  INVX0 U1 ( .INP(B[1]), .ZN(n8) );
  NAND2X1 U2 ( .IN1(n1), .IN2(B[0]), .QN(carry[1]) );
  INVX0 U3 ( .INP(A[0]), .ZN(n1) );
  INVX0 U4 ( .INP(B[2]), .ZN(n7) );
  INVX0 U5 ( .INP(B[3]), .ZN(n6) );
  INVX0 U6 ( .INP(B[4]), .ZN(n5) );
  INVX0 U7 ( .INP(B[5]), .ZN(n4) );
  INVX0 U8 ( .INP(B[6]), .ZN(n3) );
  INVX0 U9 ( .INP(B[7]), .ZN(n2) );
  XOR2X1 U10 ( .IN1(B[0]), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module combined_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[8]), .IN2(carry[8]), .Q(SUM[8]) );
  XOR2X1 U3 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module combined_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;
  assign SUM[23] = carry[23];

  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module combined ( clk, reset, exponent_a, exponent_b, fraction_a, fraction_b, 
        sign_a, sign_b, new_sign_o, new_exponent_o, combined_a_o, combined_b_o, 
        combined_negative_b_o, add_exponent_a, add_exponent_b, 
        add_difference_o, add_zero_flag_o, add_greater_flag_o, 
        add_lesser_flag_o, add_sign_a, add_sign_b, add_sign_a2, add_sign_b2, 
        add_fraction_a, add_fraction_b, add_fraction_a2, add_fraction_b2, 
        add_exponent_a2, s, s2 );
  input [7:0] exponent_a;
  input [7:0] exponent_b;
  input [22:0] fraction_a;
  input [22:0] fraction_b;
  output [8:0] new_exponent_o;
  output [24:0] combined_a_o;
  output [24:0] combined_b_o;
  output [24:0] combined_negative_b_o;
  input [7:0] add_exponent_a;
  input [7:0] add_exponent_b;
  output [7:0] add_difference_o;
  input [22:0] add_fraction_a;
  input [22:0] add_fraction_b;
  output [22:0] add_fraction_a2;
  output [22:0] add_fraction_b2;
  output [7:0] add_exponent_a2;
  input clk, reset, sign_a, sign_b, add_sign_a, add_sign_b, s;
  output new_sign_o, add_zero_flag_o, add_greater_flag_o, add_lesser_flag_o,
         add_sign_a2, add_sign_b2, s2;
  wire   new_sign, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         add_greater_flag, add_lesser_flag, N48, N49, N50, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, N9, N8, N7, N6, N5, N12, N11, N10, N45,
         N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31,
         N30, N29, N28, N27, N26, N25, N24, N23,
         \sub_1_root_sub_0_root_sub_82/carry[2] ,
         \sub_1_root_sub_0_root_sub_82/carry[3] ,
         \sub_1_root_sub_0_root_sub_82/carry[4] ,
         \sub_1_root_sub_0_root_sub_82/carry[5] ,
         \sub_1_root_sub_0_root_sub_82/carry[6] ,
         \sub_1_root_sub_0_root_sub_82/carry[7] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79;
  wire   [8:0] new_exponent;
  wire   [24:0] combined_negative_b;
  wire   [7:0] add_difference;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFFARX1 \combined_negative_b_o_reg[24]  ( .D(1'b1), .CLK(clk), .RSTB(n17), 
        .Q(combined_negative_b_o[24]) );
  DFFARX1 \combined_negative_b_o_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[23]) );
  DFFARX1 \combined_negative_b_o_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[22]) );
  DFFARX1 \combined_negative_b_o_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[21]) );
  DFFARX1 \combined_negative_b_o_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[20]) );
  DFFARX1 \combined_negative_b_o_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[19]) );
  DFFARX1 \combined_negative_b_o_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n17), .Q(combined_negative_b_o[18]) );
  DFFARX1 \combined_negative_b_o_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[17]) );
  DFFARX1 \combined_negative_b_o_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[16]) );
  DFFARX1 \combined_negative_b_o_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[15]) );
  DFFARX1 \combined_negative_b_o_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[14]) );
  DFFARX1 \combined_negative_b_o_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[13]) );
  DFFARX1 \combined_negative_b_o_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[12]) );
  DFFARX1 \combined_negative_b_o_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[11]) );
  DFFARX1 \combined_negative_b_o_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[10]) );
  DFFARX1 \combined_negative_b_o_reg[9]  ( .D(combined_negative_b[9]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[9]) );
  DFFARX1 \combined_negative_b_o_reg[8]  ( .D(combined_negative_b[8]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[8]) );
  DFFARX1 \combined_negative_b_o_reg[7]  ( .D(combined_negative_b[7]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[7]) );
  DFFARX1 \combined_negative_b_o_reg[6]  ( .D(combined_negative_b[6]), .CLK(
        clk), .RSTB(n16), .Q(combined_negative_b_o[6]) );
  DFFARX1 \combined_negative_b_o_reg[5]  ( .D(combined_negative_b[5]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[5]) );
  DFFARX1 \combined_negative_b_o_reg[4]  ( .D(combined_negative_b[4]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[4]) );
  DFFARX1 \combined_negative_b_o_reg[3]  ( .D(combined_negative_b[3]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[3]) );
  DFFARX1 \combined_negative_b_o_reg[2]  ( .D(combined_negative_b[2]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[2]) );
  DFFARX1 \combined_negative_b_o_reg[1]  ( .D(combined_negative_b[1]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[1]) );
  DFFARX1 \combined_negative_b_o_reg[0]  ( .D(combined_negative_b[0]), .CLK(
        clk), .RSTB(n15), .Q(combined_negative_b_o[0]) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n15), .Q(s2) );
  DFFARX1 new_sign_o_reg ( .D(new_sign), .CLK(clk), .RSTB(n15), .Q(new_sign_o)
         );
  DFFARX1 \new_exponent_o_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n15), 
        .Q(new_exponent_o[8]) );
  DFFARX1 \new_exponent_o_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n15), 
        .Q(new_exponent_o[7]) );
  DFFARX1 \new_exponent_o_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n15), 
        .Q(new_exponent_o[6]) );
  DFFARX1 \new_exponent_o_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n15), 
        .Q(new_exponent_o[5]) );
  DFFARX1 \new_exponent_o_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n14), 
        .Q(new_exponent_o[4]) );
  DFFARX1 \new_exponent_o_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n14), 
        .Q(new_exponent_o[3]) );
  DFFARX1 \new_exponent_o_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n14), 
        .Q(new_exponent_o[2]) );
  DFFARX1 \new_exponent_o_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n14), 
        .Q(new_exponent_o[1]) );
  DFFARX1 \new_exponent_o_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n14), 
        .Q(new_exponent_o[0]) );
  DFFARX1 \combined_a_o_reg[23]  ( .D(1'b1), .CLK(clk), .RSTB(n14), .Q(
        combined_a_o[23]) );
  DFFARX1 \combined_a_o_reg[22]  ( .D(fraction_a[22]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[22]) );
  DFFARX1 \combined_a_o_reg[21]  ( .D(fraction_a[21]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[21]) );
  DFFARX1 \combined_a_o_reg[20]  ( .D(fraction_a[20]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[20]) );
  DFFARX1 \combined_a_o_reg[19]  ( .D(fraction_a[19]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[19]) );
  DFFARX1 \combined_a_o_reg[18]  ( .D(fraction_a[18]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[18]) );
  DFFARX1 \combined_a_o_reg[17]  ( .D(fraction_a[17]), .CLK(clk), .RSTB(n14), 
        .Q(combined_a_o[17]) );
  DFFARX1 \combined_a_o_reg[16]  ( .D(fraction_a[16]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[16]) );
  DFFARX1 \combined_a_o_reg[15]  ( .D(fraction_a[15]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[15]) );
  DFFARX1 \combined_a_o_reg[14]  ( .D(fraction_a[14]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[14]) );
  DFFARX1 \combined_a_o_reg[13]  ( .D(fraction_a[13]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[13]) );
  DFFARX1 \combined_a_o_reg[12]  ( .D(fraction_a[12]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[12]) );
  DFFARX1 \combined_a_o_reg[11]  ( .D(fraction_a[11]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[11]) );
  DFFARX1 \combined_a_o_reg[10]  ( .D(fraction_a[10]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[10]) );
  DFFARX1 \combined_a_o_reg[9]  ( .D(fraction_a[9]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[9]) );
  DFFARX1 \combined_a_o_reg[8]  ( .D(fraction_a[8]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[8]) );
  DFFARX1 \combined_a_o_reg[7]  ( .D(fraction_a[7]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[7]) );
  DFFARX1 \combined_a_o_reg[6]  ( .D(fraction_a[6]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[6]) );
  DFFARX1 \combined_a_o_reg[5]  ( .D(fraction_a[5]), .CLK(clk), .RSTB(n13), 
        .Q(combined_a_o[5]) );
  DFFARX1 \combined_a_o_reg[4]  ( .D(fraction_a[4]), .CLK(clk), .RSTB(n12), 
        .Q(combined_a_o[4]) );
  DFFARX1 \combined_a_o_reg[3]  ( .D(fraction_a[3]), .CLK(clk), .RSTB(n12), 
        .Q(combined_a_o[3]) );
  DFFARX1 \combined_a_o_reg[2]  ( .D(fraction_a[2]), .CLK(clk), .RSTB(n12), 
        .Q(combined_a_o[2]) );
  DFFARX1 \combined_a_o_reg[1]  ( .D(fraction_a[1]), .CLK(clk), .RSTB(n12), 
        .Q(combined_a_o[1]) );
  DFFARX1 \combined_a_o_reg[0]  ( .D(fraction_a[0]), .CLK(clk), .RSTB(n12), 
        .Q(combined_a_o[0]) );
  DFFARX1 \combined_b_o_reg[23]  ( .D(1'b1), .CLK(clk), .RSTB(n12), .Q(
        combined_b_o[23]) );
  DFFARX1 \combined_b_o_reg[22]  ( .D(fraction_b[22]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[22]) );
  DFFARX1 \combined_b_o_reg[21]  ( .D(fraction_b[21]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[21]) );
  DFFARX1 \combined_b_o_reg[20]  ( .D(fraction_b[20]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[20]) );
  DFFARX1 \combined_b_o_reg[19]  ( .D(fraction_b[19]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[19]) );
  DFFARX1 \combined_b_o_reg[18]  ( .D(fraction_b[18]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[18]) );
  DFFARX1 \combined_b_o_reg[17]  ( .D(fraction_b[17]), .CLK(clk), .RSTB(n12), 
        .Q(combined_b_o[17]) );
  DFFARX1 \combined_b_o_reg[16]  ( .D(fraction_b[16]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[16]) );
  DFFARX1 \combined_b_o_reg[15]  ( .D(fraction_b[15]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[15]) );
  DFFARX1 \combined_b_o_reg[14]  ( .D(fraction_b[14]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[14]) );
  DFFARX1 \combined_b_o_reg[13]  ( .D(fraction_b[13]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[13]) );
  DFFARX1 \combined_b_o_reg[12]  ( .D(fraction_b[12]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[12]) );
  DFFARX1 \combined_b_o_reg[11]  ( .D(fraction_b[11]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[11]) );
  DFFARX1 \combined_b_o_reg[10]  ( .D(fraction_b[10]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[10]) );
  DFFARX1 \combined_b_o_reg[9]  ( .D(fraction_b[9]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[9]) );
  DFFARX1 \combined_b_o_reg[8]  ( .D(fraction_b[8]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[8]) );
  DFFARX1 \combined_b_o_reg[7]  ( .D(fraction_b[7]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[7]) );
  DFFARX1 \combined_b_o_reg[6]  ( .D(fraction_b[6]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[6]) );
  DFFARX1 \combined_b_o_reg[5]  ( .D(fraction_b[5]), .CLK(clk), .RSTB(n11), 
        .Q(combined_b_o[5]) );
  DFFARX1 \combined_b_o_reg[4]  ( .D(fraction_b[4]), .CLK(clk), .RSTB(n10), 
        .Q(combined_b_o[4]) );
  DFFARX1 \combined_b_o_reg[3]  ( .D(fraction_b[3]), .CLK(clk), .RSTB(n10), 
        .Q(combined_b_o[3]) );
  DFFARX1 \combined_b_o_reg[2]  ( .D(fraction_b[2]), .CLK(clk), .RSTB(n10), 
        .Q(combined_b_o[2]) );
  DFFARX1 \combined_b_o_reg[1]  ( .D(fraction_b[1]), .CLK(clk), .RSTB(n10), 
        .Q(combined_b_o[1]) );
  DFFARX1 \combined_b_o_reg[0]  ( .D(fraction_b[0]), .CLK(clk), .RSTB(n10), 
        .Q(combined_b_o[0]) );
  DFFARX1 add_sign_b2_reg ( .D(add_sign_b), .CLK(clk), .RSTB(n10), .Q(
        add_sign_b2) );
  DFFARX1 \add_exponent_a2_reg[7]  ( .D(add_exponent_a[7]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[7]) );
  DFFARX1 \add_exponent_a2_reg[6]  ( .D(add_exponent_a[6]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[6]) );
  DFFARX1 \add_exponent_a2_reg[5]  ( .D(add_exponent_a[5]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[5]) );
  DFFARX1 \add_exponent_a2_reg[4]  ( .D(add_exponent_a[4]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[4]) );
  DFFARX1 \add_exponent_a2_reg[3]  ( .D(add_exponent_a[3]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[3]) );
  DFFARX1 \add_exponent_a2_reg[2]  ( .D(add_exponent_a[2]), .CLK(clk), .RSTB(
        n10), .Q(add_exponent_a2[2]) );
  DFFARX1 \add_exponent_a2_reg[1]  ( .D(add_exponent_a[1]), .CLK(clk), .RSTB(
        n9), .Q(add_exponent_a2[1]) );
  DFFARX1 \add_exponent_a2_reg[0]  ( .D(add_exponent_a[0]), .CLK(clk), .RSTB(
        n9), .Q(add_exponent_a2[0]) );
  DFFARX1 \add_difference_o_reg[7]  ( .D(add_difference[7]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[7]) );
  DFFARX1 \add_difference_o_reg[6]  ( .D(add_difference[6]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[6]) );
  DFFARX1 \add_difference_o_reg[5]  ( .D(add_difference[5]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[5]) );
  DFFARX1 \add_difference_o_reg[4]  ( .D(add_difference[4]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[4]) );
  DFFARX1 \add_difference_o_reg[3]  ( .D(add_difference[3]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[3]) );
  DFFARX1 \add_difference_o_reg[2]  ( .D(add_difference[2]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[2]) );
  DFFARX1 \add_difference_o_reg[1]  ( .D(add_difference[1]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[1]) );
  DFFARX1 \add_difference_o_reg[0]  ( .D(add_difference[0]), .CLK(clk), .RSTB(
        n9), .Q(add_difference_o[0]) );
  DFFARX1 add_zero_flag_o_reg ( .D(N48), .CLK(clk), .RSTB(n9), .Q(
        add_zero_flag_o) );
  DFFARX1 add_greater_flag_o_reg ( .D(add_greater_flag), .CLK(clk), .RSTB(n9), 
        .Q(add_greater_flag_o) );
  DFFARX1 add_lesser_flag_o_reg ( .D(add_lesser_flag), .CLK(clk), .RSTB(n8), 
        .Q(add_lesser_flag_o) );
  DFFARX1 \add_fraction_a2_reg[22]  ( .D(add_fraction_a[22]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[22]) );
  DFFARX1 \add_fraction_a2_reg[21]  ( .D(add_fraction_a[21]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[21]) );
  DFFARX1 \add_fraction_a2_reg[20]  ( .D(add_fraction_a[20]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[20]) );
  DFFARX1 \add_fraction_a2_reg[19]  ( .D(add_fraction_a[19]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[19]) );
  DFFARX1 \add_fraction_a2_reg[18]  ( .D(add_fraction_a[18]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[18]) );
  DFFARX1 \add_fraction_a2_reg[17]  ( .D(add_fraction_a[17]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[17]) );
  DFFARX1 \add_fraction_a2_reg[16]  ( .D(add_fraction_a[16]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[16]) );
  DFFARX1 \add_fraction_a2_reg[15]  ( .D(add_fraction_a[15]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[15]) );
  DFFARX1 \add_fraction_a2_reg[14]  ( .D(add_fraction_a[14]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[14]) );
  DFFARX1 \add_fraction_a2_reg[13]  ( .D(add_fraction_a[13]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[13]) );
  DFFARX1 \add_fraction_a2_reg[12]  ( .D(add_fraction_a[12]), .CLK(clk), 
        .RSTB(n8), .Q(add_fraction_a2[12]) );
  DFFARX1 \add_fraction_a2_reg[11]  ( .D(add_fraction_a[11]), .CLK(clk), 
        .RSTB(n7), .Q(add_fraction_a2[11]) );
  DFFARX1 \add_fraction_a2_reg[10]  ( .D(add_fraction_a[10]), .CLK(clk), 
        .RSTB(n7), .Q(add_fraction_a2[10]) );
  DFFARX1 \add_fraction_a2_reg[9]  ( .D(add_fraction_a[9]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[9]) );
  DFFARX1 \add_fraction_a2_reg[8]  ( .D(add_fraction_a[8]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[8]) );
  DFFARX1 \add_fraction_a2_reg[7]  ( .D(add_fraction_a[7]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[7]) );
  DFFARX1 \add_fraction_a2_reg[6]  ( .D(add_fraction_a[6]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[6]) );
  DFFARX1 \add_fraction_a2_reg[5]  ( .D(add_fraction_a[5]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[5]) );
  DFFARX1 \add_fraction_a2_reg[4]  ( .D(add_fraction_a[4]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[4]) );
  DFFARX1 \add_fraction_a2_reg[3]  ( .D(add_fraction_a[3]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[3]) );
  DFFARX1 \add_fraction_a2_reg[2]  ( .D(add_fraction_a[2]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[2]) );
  DFFARX1 \add_fraction_a2_reg[1]  ( .D(add_fraction_a[1]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[1]) );
  DFFARX1 \add_fraction_a2_reg[0]  ( .D(add_fraction_a[0]), .CLK(clk), .RSTB(
        n7), .Q(add_fraction_a2[0]) );
  DFFARX1 \add_fraction_b2_reg[22]  ( .D(add_fraction_b[22]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[22]) );
  DFFARX1 \add_fraction_b2_reg[21]  ( .D(add_fraction_b[21]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[21]) );
  DFFARX1 \add_fraction_b2_reg[20]  ( .D(add_fraction_b[20]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[20]) );
  DFFARX1 \add_fraction_b2_reg[19]  ( .D(add_fraction_b[19]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[19]) );
  DFFARX1 \add_fraction_b2_reg[18]  ( .D(add_fraction_b[18]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[18]) );
  DFFARX1 \add_fraction_b2_reg[17]  ( .D(add_fraction_b[17]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[17]) );
  DFFARX1 \add_fraction_b2_reg[16]  ( .D(add_fraction_b[16]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[16]) );
  DFFARX1 \add_fraction_b2_reg[15]  ( .D(add_fraction_b[15]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[15]) );
  DFFARX1 \add_fraction_b2_reg[14]  ( .D(add_fraction_b[14]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[14]) );
  DFFARX1 \add_fraction_b2_reg[13]  ( .D(add_fraction_b[13]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[13]) );
  DFFARX1 \add_fraction_b2_reg[12]  ( .D(add_fraction_b[12]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[12]) );
  DFFARX1 \add_fraction_b2_reg[11]  ( .D(add_fraction_b[11]), .CLK(clk), 
        .RSTB(n6), .Q(add_fraction_b2[11]) );
  DFFARX1 \add_fraction_b2_reg[10]  ( .D(add_fraction_b[10]), .CLK(clk), 
        .RSTB(n5), .Q(add_fraction_b2[10]) );
  DFFARX1 \add_fraction_b2_reg[9]  ( .D(add_fraction_b[9]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[9]) );
  DFFARX1 \add_fraction_b2_reg[8]  ( .D(add_fraction_b[8]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[8]) );
  DFFARX1 \add_fraction_b2_reg[7]  ( .D(add_fraction_b[7]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[7]) );
  DFFARX1 \add_fraction_b2_reg[6]  ( .D(add_fraction_b[6]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[6]) );
  DFFARX1 \add_fraction_b2_reg[5]  ( .D(add_fraction_b[5]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[5]) );
  DFFARX1 \add_fraction_b2_reg[4]  ( .D(add_fraction_b[4]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[4]) );
  DFFARX1 \add_fraction_b2_reg[3]  ( .D(add_fraction_b[3]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[3]) );
  DFFARX1 \add_fraction_b2_reg[2]  ( .D(add_fraction_b[2]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[2]) );
  DFFARX1 \add_fraction_b2_reg[1]  ( .D(add_fraction_b[1]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[1]) );
  DFFARX1 \add_fraction_b2_reg[0]  ( .D(add_fraction_b[0]), .CLK(clk), .RSTB(
        n5), .Q(add_fraction_b2[0]) );
  DFFARX1 add_sign_a2_reg ( .D(add_sign_a), .CLK(clk), .RSTB(n5), .Q(
        add_sign_a2) );
  XOR2X1 U11 ( .IN1(sign_b), .IN2(sign_a), .Q(new_sign) );
  AND2X1 U12 ( .IN1(N22), .IN2(n21), .Q(new_exponent[8]) );
  AND2X1 U13 ( .IN1(N21), .IN2(n21), .Q(new_exponent[7]) );
  AND2X1 U14 ( .IN1(N20), .IN2(n21), .Q(new_exponent[6]) );
  AND2X1 U15 ( .IN1(N19), .IN2(n21), .Q(new_exponent[5]) );
  AND2X1 U16 ( .IN1(N18), .IN2(n21), .Q(new_exponent[4]) );
  AND2X1 U17 ( .IN1(N17), .IN2(n21), .Q(new_exponent[3]) );
  AND2X1 U18 ( .IN1(N16), .IN2(n21), .Q(new_exponent[2]) );
  AND2X1 U19 ( .IN1(N15), .IN2(n21), .Q(new_exponent[1]) );
  AND2X1 U20 ( .IN1(N14), .IN2(n21), .Q(new_exponent[0]) );
  NAND4X0 U22 ( .IN1(n26), .IN2(n27), .IN3(n28), .IN4(n29), .QN(n25) );
  NOR4X0 U23 ( .IN1(fraction_b[15]), .IN2(fraction_b[14]), .IN3(fraction_b[13]), .IN4(fraction_b[12]), .QN(n29) );
  NOR4X0 U24 ( .IN1(fraction_b[11]), .IN2(fraction_b[10]), .IN3(fraction_b[0]), 
        .IN4(fraction_a[9]), .QN(n28) );
  NOR4X0 U25 ( .IN1(fraction_a[8]), .IN2(fraction_a[7]), .IN3(fraction_a[6]), 
        .IN4(fraction_a[5]), .QN(n27) );
  NOR3X0 U26 ( .IN1(fraction_a[2]), .IN2(fraction_a[4]), .IN3(fraction_a[3]), 
        .QN(n26) );
  NAND4X0 U27 ( .IN1(n30), .IN2(n31), .IN3(n32), .IN4(n33), .QN(n24) );
  NOR4X0 U28 ( .IN1(fraction_b[9]), .IN2(fraction_b[8]), .IN3(fraction_b[7]), 
        .IN4(fraction_b[6]), .QN(n33) );
  NOR4X0 U29 ( .IN1(fraction_b[5]), .IN2(fraction_b[4]), .IN3(fraction_b[3]), 
        .IN4(fraction_b[2]), .QN(n32) );
  NOR4X0 U30 ( .IN1(fraction_b[22]), .IN2(fraction_b[21]), .IN3(fraction_b[20]), .IN4(fraction_b[1]), .QN(n31) );
  NOR4X0 U31 ( .IN1(fraction_b[19]), .IN2(fraction_b[18]), .IN3(fraction_b[17]), .IN4(fraction_b[16]), .QN(n30) );
  NAND4X0 U32 ( .IN1(n34), .IN2(n35), .IN3(n36), .IN4(n37), .QN(n23) );
  NOR4X0 U33 ( .IN1(exponent_b[6]), .IN2(exponent_b[5]), .IN3(exponent_b[4]), 
        .IN4(exponent_b[3]), .QN(n37) );
  NOR4X0 U34 ( .IN1(exponent_b[2]), .IN2(exponent_b[1]), .IN3(exponent_b[0]), 
        .IN4(exponent_a[7]), .QN(n36) );
  NOR4X0 U35 ( .IN1(exponent_a[6]), .IN2(exponent_a[5]), .IN3(exponent_a[4]), 
        .IN4(exponent_a[3]), .QN(n35) );
  NOR3X0 U36 ( .IN1(exponent_a[0]), .IN2(exponent_a[2]), .IN3(exponent_a[1]), 
        .QN(n34) );
  NAND4X0 U37 ( .IN1(n38), .IN2(n39), .IN3(n40), .IN4(n41), .QN(n22) );
  NOR4X0 U38 ( .IN1(fraction_a[22]), .IN2(fraction_a[21]), .IN3(fraction_a[20]), .IN4(fraction_a[1]), .QN(n41) );
  NOR4X0 U39 ( .IN1(fraction_a[19]), .IN2(fraction_a[18]), .IN3(fraction_a[17]), .IN4(fraction_a[16]), .QN(n40) );
  NOR4X0 U40 ( .IN1(fraction_a[15]), .IN2(fraction_a[14]), .IN3(fraction_a[13]), .IN4(fraction_a[12]), .QN(n39) );
  NOR4X0 U41 ( .IN1(fraction_a[11]), .IN2(fraction_a[10]), .IN3(fraction_a[0]), 
        .IN4(exponent_b[7]), .QN(n38) );
  AND2X1 U42 ( .IN1(N50), .IN2(n42), .Q(add_lesser_flag) );
  AO22X1 U43 ( .IN1(N64), .IN2(add_greater_flag), .IN3(N72), .IN4(n42), .Q(
        add_difference[7]) );
  AO22X1 U44 ( .IN1(N63), .IN2(add_greater_flag), .IN3(N71), .IN4(n42), .Q(
        add_difference[6]) );
  AO22X1 U45 ( .IN1(N62), .IN2(add_greater_flag), .IN3(N70), .IN4(n42), .Q(
        add_difference[5]) );
  AO22X1 U46 ( .IN1(N61), .IN2(add_greater_flag), .IN3(N69), .IN4(n42), .Q(
        add_difference[4]) );
  AO22X1 U47 ( .IN1(N60), .IN2(add_greater_flag), .IN3(N68), .IN4(n42), .Q(
        add_difference[3]) );
  AO22X1 U48 ( .IN1(N59), .IN2(add_greater_flag), .IN3(N67), .IN4(n42), .Q(
        add_difference[2]) );
  AO22X1 U49 ( .IN1(N58), .IN2(add_greater_flag), .IN3(N66), .IN4(n42), .Q(
        add_difference[1]) );
  AO22X1 U50 ( .IN1(N57), .IN2(add_greater_flag), .IN3(N65), .IN4(n42), .Q(
        add_difference[0]) );
  combined_DW01_sub_0 sub_165 ( .A(add_exponent_b), .B(add_exponent_a), .CI(
        1'b0), .DIFF({N72, N71, N70, N69, N68, N67, N66, N65}) );
  combined_DW01_sub_1 sub_163 ( .A(add_exponent_a), .B(add_exponent_b), .CI(
        1'b0), .DIFF({N64, N63, N62, N61, N60, N59, N58, N57}) );
  combined_DW01_add_0 add_0_root_sub_0_root_sub_82 ( .A({1'b0, exponent_b}), 
        .B({n3, N12, N11, N10, N9, N8, N7, N6, N5}), .CI(1'b0), .SUM({N22, N21, 
        N20, N19, N18, N17, N16, N15, N14}) );
  combined_DW01_inc_0 add_91 ( .A({1'b1, 1'b0, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23}), .SUM({SYNOPSYS_UNCONNECTED__0, 
        combined_negative_b[23:0]}) );
  NOR2X0 U3 ( .IN1(exponent_a[7]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[7] ), .QN(n3) );
  NBUFFX2 U4 ( .INP(n4), .Z(n5) );
  NBUFFX2 U5 ( .INP(n4), .Z(n6) );
  NBUFFX2 U8 ( .INP(n4), .Z(n7) );
  NBUFFX2 U9 ( .INP(n4), .Z(n8) );
  NBUFFX2 U10 ( .INP(n4), .Z(n9) );
  NBUFFX2 U21 ( .INP(n4), .Z(n10) );
  NBUFFX2 U51 ( .INP(n4), .Z(n11) );
  NBUFFX2 U52 ( .INP(n4), .Z(n12) );
  NBUFFX2 U53 ( .INP(n4), .Z(n13) );
  NBUFFX2 U54 ( .INP(n4), .Z(n14) );
  NBUFFX2 U55 ( .INP(n4), .Z(n15) );
  NBUFFX2 U56 ( .INP(n4), .Z(n16) );
  NBUFFX2 U57 ( .INP(n4), .Z(n17) );
  NOR2X0 U58 ( .IN1(N48), .IN2(N49), .QN(n42) );
  NOR2X0 U59 ( .IN1(n79), .IN2(N48), .QN(add_greater_flag) );
  INVX0 U60 ( .INP(N49), .ZN(n79) );
  INVX0 U61 ( .INP(n18), .ZN(n74) );
  OR4X1 U62 ( .IN1(n22), .IN2(n23), .IN3(n24), .IN4(n25), .Q(n21) );
  NBUFFX2 U63 ( .INP(reset), .Z(n4) );
  INVX0 U64 ( .INP(fraction_b[1]), .ZN(N24) );
  INVX0 U65 ( .INP(fraction_b[2]), .ZN(N25) );
  INVX0 U66 ( .INP(fraction_b[3]), .ZN(N26) );
  INVX0 U67 ( .INP(fraction_b[4]), .ZN(N27) );
  INVX0 U68 ( .INP(fraction_b[5]), .ZN(N28) );
  INVX0 U69 ( .INP(fraction_b[6]), .ZN(N29) );
  INVX0 U70 ( .INP(fraction_b[7]), .ZN(N30) );
  INVX0 U71 ( .INP(fraction_b[8]), .ZN(N31) );
  INVX0 U72 ( .INP(fraction_b[9]), .ZN(N32) );
  INVX0 U73 ( .INP(fraction_b[10]), .ZN(N33) );
  INVX0 U74 ( .INP(fraction_b[11]), .ZN(N34) );
  INVX0 U75 ( .INP(fraction_b[12]), .ZN(N35) );
  INVX0 U76 ( .INP(fraction_b[13]), .ZN(N36) );
  INVX0 U77 ( .INP(fraction_b[14]), .ZN(N37) );
  INVX0 U78 ( .INP(fraction_b[15]), .ZN(N38) );
  INVX0 U79 ( .INP(fraction_b[16]), .ZN(N39) );
  INVX0 U80 ( .INP(fraction_b[17]), .ZN(N40) );
  INVX0 U81 ( .INP(fraction_b[18]), .ZN(N41) );
  INVX0 U82 ( .INP(fraction_b[19]), .ZN(N42) );
  INVX0 U83 ( .INP(fraction_b[20]), .ZN(N43) );
  INVX0 U84 ( .INP(fraction_b[21]), .ZN(N44) );
  INVX0 U85 ( .INP(fraction_b[22]), .ZN(N45) );
  INVX0 U86 ( .INP(fraction_b[0]), .ZN(N23) );
  INVX0 U87 ( .INP(exponent_a[0]), .ZN(N5) );
  INVX0 U88 ( .INP(add_exponent_b[1]), .ZN(n70) );
  INVX0 U89 ( .INP(add_exponent_a[1]), .ZN(n75) );
  INVX0 U90 ( .INP(add_exponent_a[2]), .ZN(n76) );
  INVX0 U91 ( .INP(add_exponent_a[4]), .ZN(n77) );
  INVX0 U92 ( .INP(add_exponent_b[0]), .ZN(n69) );
  INVX0 U93 ( .INP(add_exponent_b[6]), .ZN(n73) );
  INVX0 U94 ( .INP(add_exponent_b[3]), .ZN(n71) );
  INVX0 U95 ( .INP(add_exponent_b[5]), .ZN(n72) );
  INVX0 U96 ( .INP(add_exponent_a[7]), .ZN(n78) );
  XNOR2X1 U97 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[7] ), .IN2(
        exponent_a[7]), .Q(N12) );
  AND2X1 U98 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[6] ), .IN2(
        exponent_a[6]), .Q(\sub_1_root_sub_0_root_sub_82/carry[7] ) );
  XOR2X1 U99 ( .IN1(exponent_a[6]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[6] ), .Q(N11) );
  AND2X1 U100 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[5] ), .IN2(
        exponent_a[5]), .Q(\sub_1_root_sub_0_root_sub_82/carry[6] ) );
  XOR2X1 U101 ( .IN1(exponent_a[5]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[5] ), .Q(N10) );
  AND2X1 U102 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[4] ), .IN2(
        exponent_a[4]), .Q(\sub_1_root_sub_0_root_sub_82/carry[5] ) );
  XOR2X1 U103 ( .IN1(exponent_a[4]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[4] ), .Q(N9) );
  AND2X1 U104 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[3] ), .IN2(
        exponent_a[3]), .Q(\sub_1_root_sub_0_root_sub_82/carry[4] ) );
  XOR2X1 U105 ( .IN1(exponent_a[3]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[3] ), .Q(N8) );
  AND2X1 U106 ( .IN1(\sub_1_root_sub_0_root_sub_82/carry[2] ), .IN2(
        exponent_a[2]), .Q(\sub_1_root_sub_0_root_sub_82/carry[3] ) );
  XOR2X1 U107 ( .IN1(exponent_a[2]), .IN2(
        \sub_1_root_sub_0_root_sub_82/carry[2] ), .Q(N7) );
  AND2X1 U108 ( .IN1(exponent_a[0]), .IN2(exponent_a[1]), .Q(
        \sub_1_root_sub_0_root_sub_82/carry[2] ) );
  XOR2X1 U109 ( .IN1(exponent_a[1]), .IN2(exponent_a[0]), .Q(N6) );
  NOR2X0 U110 ( .IN1(n78), .IN2(add_exponent_b[7]), .QN(n66) );
  NOR2X0 U111 ( .IN1(n69), .IN2(add_exponent_a[0]), .QN(n18) );
  NAND2X0 U112 ( .IN1(n18), .IN2(n75), .QN(n19) );
  OR2X1 U113 ( .IN1(n76), .IN2(add_exponent_b[2]), .Q(n54) );
  NAND2X0 U114 ( .IN1(add_exponent_b[2]), .IN2(n76), .QN(n20) );
  NAND2X0 U115 ( .IN1(n54), .IN2(n20), .QN(n50) );
  AO221X1 U116 ( .IN1(n19), .IN2(n70), .IN3(add_exponent_a[1]), .IN4(n74), 
        .IN5(n50), .Q(n43) );
  OR2X1 U117 ( .IN1(n71), .IN2(add_exponent_a[3]), .Q(n57) );
  NAND3X0 U118 ( .IN1(n43), .IN2(n20), .IN3(n57), .QN(n44) );
  NAND2X0 U119 ( .IN1(add_exponent_a[3]), .IN2(n71), .QN(n55) );
  OR2X1 U120 ( .IN1(n77), .IN2(add_exponent_b[4]), .Q(n60) );
  NAND2X0 U121 ( .IN1(add_exponent_b[4]), .IN2(n77), .QN(n45) );
  AND2X1 U122 ( .IN1(n60), .IN2(n45), .Q(n56) );
  NAND3X0 U123 ( .IN1(n44), .IN2(n55), .IN3(n56), .QN(n46) );
  OR2X1 U124 ( .IN1(n72), .IN2(add_exponent_a[5]), .Q(n63) );
  NAND3X0 U125 ( .IN1(n46), .IN2(n45), .IN3(n63), .QN(n47) );
  NAND2X0 U126 ( .IN1(add_exponent_a[5]), .IN2(n72), .QN(n61) );
  XOR2X1 U127 ( .IN1(add_exponent_a[6]), .IN2(n73), .Q(n62) );
  NAND3X0 U128 ( .IN1(n47), .IN2(n61), .IN3(n62), .QN(n48) );
  OA21X1 U129 ( .IN1(add_exponent_a[6]), .IN2(n73), .IN3(n48), .Q(n49) );
  NAND2X0 U130 ( .IN1(add_exponent_b[7]), .IN2(n78), .QN(n68) );
  OAI21X1 U131 ( .IN1(n66), .IN2(n49), .IN3(n68), .QN(N50) );
  NAND2X0 U132 ( .IN1(add_exponent_a[0]), .IN2(n69), .QN(n51) );
  OR2X1 U133 ( .IN1(n51), .IN2(n75), .Q(n52) );
  AO221X1 U134 ( .IN1(add_exponent_b[1]), .IN2(n52), .IN3(n51), .IN4(n75), 
        .IN5(n50), .Q(n53) );
  NAND3X0 U135 ( .IN1(n55), .IN2(n54), .IN3(n53), .QN(n58) );
  NAND3X0 U136 ( .IN1(n58), .IN2(n57), .IN3(n56), .QN(n59) );
  NAND3X0 U137 ( .IN1(n61), .IN2(n60), .IN3(n59), .QN(n64) );
  AND3X1 U138 ( .IN1(n64), .IN2(n63), .IN3(n62), .Q(n65) );
  AO21X1 U139 ( .IN1(n73), .IN2(add_exponent_a[6]), .IN3(n65), .Q(n67) );
  AO21X1 U140 ( .IN1(n68), .IN2(n67), .IN3(n66), .Q(N49) );
  NOR2X0 U141 ( .IN1(N50), .IN2(N49), .QN(N48) );
endmodule


module booth_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .IN1(A[7]), .IN2(B[7]), .IN3(carry[7]), .Q(SUM[7]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module booth_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND3X0 U3 ( .IN1(n65), .IN2(n66), .IN3(n1), .QN(n69) );
  AO221X1 U4 ( .IN1(A[21]), .IN2(SH[0]), .IN3(A[22]), .IN4(SH[1]), .IN5(n102), 
        .Q(n49) );
  INVX0 U5 ( .INP(n55), .ZN(n10) );
  INVX0 U6 ( .INP(n68), .ZN(n7) );
  INVX0 U7 ( .INP(n75), .ZN(n4) );
  INVX0 U8 ( .INP(n80), .ZN(n5) );
  INVX0 U9 ( .INP(n82), .ZN(n6) );
  INVX0 U10 ( .INP(n91), .ZN(n3) );
  INVX0 U11 ( .INP(n56), .ZN(n9) );
  INVX0 U12 ( .INP(n78), .ZN(n12) );
  AND2X1 U13 ( .IN1(n21), .IN2(SH[2]), .Q(n31) );
  MUX21X1 U14 ( .IN1(n40), .IN2(n84), .S(SH[2]), .Q(n82) );
  MUX21X1 U15 ( .IN1(n32), .IN2(n10), .S(SH[2]), .Q(n80) );
  INVX0 U16 ( .INP(n79), .ZN(n13) );
  INVX0 U17 ( .INP(n66), .ZN(n2) );
  INVX0 U18 ( .INP(SH[7]), .ZN(n1) );
  INVX0 U19 ( .INP(SH[0]), .ZN(n14) );
  INVX0 U20 ( .INP(SH[1]), .ZN(n11) );
  INVX0 U21 ( .INP(A[1]), .ZN(n18) );
  INVX0 U22 ( .INP(A[3]), .ZN(n16) );
  INVX0 U23 ( .INP(A[2]), .ZN(n17) );
  INVX0 U24 ( .INP(A[4]), .ZN(n15) );
  INVX0 U25 ( .INP(SH[2]), .ZN(n8) );
  AO222X1 U26 ( .IN1(n19), .IN2(n20), .IN3(n21), .IN4(n22), .IN5(n23), .IN6(
        n24), .Q(B[9]) );
  AO222X1 U27 ( .IN1(n19), .IN2(n25), .IN3(n21), .IN4(n26), .IN5(n23), .IN6(
        n27), .Q(B[8]) );
  AO221X1 U28 ( .IN1(n19), .IN2(n28), .IN3(n23), .IN4(n29), .IN5(n30), .Q(B[7]) );
  AO222X1 U29 ( .IN1(n31), .IN2(n32), .IN3(n33), .IN4(n10), .IN5(n34), .IN6(
        n35), .Q(n30) );
  AO221X1 U30 ( .IN1(n19), .IN2(n36), .IN3(n23), .IN4(n37), .IN5(n38), .Q(B[6]) );
  AO222X1 U31 ( .IN1(n34), .IN2(n39), .IN3(n31), .IN4(n40), .IN5(n7), .IN6(n41), .Q(n38) );
  AO221X1 U32 ( .IN1(n19), .IN2(n42), .IN3(n23), .IN4(n20), .IN5(n43), .Q(B[5]) );
  AO222X1 U33 ( .IN1(n31), .IN2(n44), .IN3(n33), .IN4(n45), .IN5(n34), .IN6(
        n24), .Q(n43) );
  AO221X1 U34 ( .IN1(n19), .IN2(n46), .IN3(n23), .IN4(n25), .IN5(n47), .Q(B[4]) );
  AO222X1 U35 ( .IN1(n31), .IN2(n48), .IN3(n33), .IN4(n49), .IN5(n34), .IN6(
        n27), .Q(n47) );
  AND2X1 U36 ( .IN1(n41), .IN2(n8), .Q(n33) );
  NOR2X0 U37 ( .IN1(n50), .IN2(SH[7]), .QN(n41) );
  NOR2X0 U38 ( .IN1(SH[7]), .IN2(n51), .QN(B[3]) );
  OA222X1 U39 ( .IN1(n52), .IN2(n2), .IN3(n5), .IN4(n50), .IN5(n53), .IN6(n54), 
        .Q(n51) );
  OA221X1 U40 ( .IN1(n55), .IN2(n16), .IN3(n56), .IN4(n15), .IN5(n57), .Q(n53)
         );
  AOI22X1 U41 ( .IN1(n12), .IN2(A[5]), .IN3(n13), .IN4(A[6]), .QN(n57) );
  AOI222X1 U42 ( .IN1(n28), .IN2(n3), .IN3(n29), .IN4(n58), .IN5(n35), .IN6(
        n59), .QN(n52) );
  AO221X1 U43 ( .IN1(A[9]), .IN2(n12), .IN3(A[10]), .IN4(n13), .IN5(n60), .Q(
        n28) );
  AO22X1 U44 ( .IN1(A[7]), .IN2(n10), .IN3(A[8]), .IN4(n9), .Q(n60) );
  NOR2X0 U45 ( .IN1(SH[7]), .IN2(n61), .QN(B[2]) );
  OA222X1 U46 ( .IN1(n62), .IN2(n2), .IN3(n6), .IN4(n50), .IN5(n63), .IN6(n54), 
        .Q(n61) );
  OA221X1 U47 ( .IN1(n55), .IN2(n17), .IN3(n56), .IN4(n16), .IN5(n64), .Q(n63)
         );
  AOI22X1 U48 ( .IN1(n12), .IN2(A[4]), .IN3(n13), .IN4(A[5]), .QN(n64) );
  NAND2X0 U49 ( .IN1(n65), .IN2(n2), .QN(n50) );
  AOI222X1 U50 ( .IN1(n36), .IN2(n3), .IN3(n37), .IN4(n58), .IN5(n39), .IN6(
        n59), .QN(n62) );
  AO221X1 U51 ( .IN1(A[8]), .IN2(n12), .IN3(A[9]), .IN4(n13), .IN5(n67), .Q(
        n36) );
  AO22X1 U52 ( .IN1(A[6]), .IN2(n10), .IN3(A[7]), .IN4(n9), .Q(n67) );
  AND2X1 U53 ( .IN1(n10), .IN2(n19), .Q(B[23]) );
  NOR2X0 U54 ( .IN1(n68), .IN2(n69), .QN(B[22]) );
  AND2X1 U55 ( .IN1(n45), .IN2(n19), .Q(B[21]) );
  AND2X1 U56 ( .IN1(n49), .IN2(n19), .Q(B[20]) );
  OA21X1 U57 ( .IN1(n70), .IN2(n71), .IN3(n1), .Q(B[1]) );
  MUX21X1 U58 ( .IN1(n4), .IN2(n72), .S(n66), .Q(n71) );
  AO222X1 U59 ( .IN1(n59), .IN2(n24), .IN3(n58), .IN4(n20), .IN5(n3), .IN6(n42), .Q(n72) );
  AO221X1 U60 ( .IN1(A[7]), .IN2(n12), .IN3(A[8]), .IN4(n13), .IN5(n73), .Q(
        n42) );
  AO22X1 U61 ( .IN1(A[5]), .IN2(n10), .IN3(A[6]), .IN4(n9), .Q(n73) );
  AO221X1 U62 ( .IN1(A[11]), .IN2(n12), .IN3(A[12]), .IN4(n13), .IN5(n74), .Q(
        n20) );
  AO22X1 U63 ( .IN1(A[9]), .IN2(n10), .IN3(A[10]), .IN4(n9), .Q(n74) );
  NOR2X0 U64 ( .IN1(n76), .IN2(n54), .QN(n70) );
  OA221X1 U65 ( .IN1(n55), .IN2(n18), .IN3(n56), .IN4(n17), .IN5(n77), .Q(n76)
         );
  OA22X1 U66 ( .IN1(n78), .IN2(n16), .IN3(n79), .IN4(n15), .Q(n77) );
  NOR2X0 U67 ( .IN1(n5), .IN2(n69), .QN(B[19]) );
  NOR2X0 U68 ( .IN1(n6), .IN2(n69), .QN(B[18]) );
  NOR2X0 U69 ( .IN1(n81), .IN2(n75), .QN(B[17]) );
  NAND2X0 U70 ( .IN1(n65), .IN2(n22), .QN(n75) );
  MUX21X1 U71 ( .IN1(n45), .IN2(n44), .S(n8), .Q(n22) );
  NOR2X0 U72 ( .IN1(n81), .IN2(n83), .QN(B[16]) );
  AO222X1 U73 ( .IN1(n19), .IN2(n35), .IN3(n34), .IN4(n10), .IN5(n23), .IN6(
        n32), .Q(B[15]) );
  AO222X1 U74 ( .IN1(n7), .IN2(n21), .IN3(n19), .IN4(n39), .IN5(n23), .IN6(n40), .Q(B[14]) );
  NAND2X0 U75 ( .IN1(n84), .IN2(n8), .QN(n68) );
  AO222X1 U76 ( .IN1(n19), .IN2(n24), .IN3(n34), .IN4(n45), .IN5(n23), .IN6(
        n44), .Q(B[13]) );
  AO221X1 U77 ( .IN1(A[19]), .IN2(n12), .IN3(A[20]), .IN4(n13), .IN5(n85), .Q(
        n44) );
  AO22X1 U78 ( .IN1(A[17]), .IN2(n10), .IN3(A[18]), .IN4(n9), .Q(n85) );
  AO221X1 U79 ( .IN1(A[22]), .IN2(n9), .IN3(A[21]), .IN4(n14), .IN5(n12), .Q(
        n45) );
  AO221X1 U80 ( .IN1(A[15]), .IN2(n12), .IN3(A[16]), .IN4(n13), .IN5(n86), .Q(
        n24) );
  AO22X1 U81 ( .IN1(A[13]), .IN2(n10), .IN3(A[14]), .IN4(n9), .Q(n86) );
  AO222X1 U82 ( .IN1(n19), .IN2(n27), .IN3(n34), .IN4(n49), .IN5(n23), .IN6(
        n48), .Q(B[12]) );
  AND2X1 U83 ( .IN1(n21), .IN2(n8), .Q(n34) );
  AO222X1 U84 ( .IN1(n21), .IN2(n80), .IN3(n19), .IN4(n29), .IN5(n23), .IN6(
        n35), .Q(B[11]) );
  AO221X1 U85 ( .IN1(A[17]), .IN2(n12), .IN3(A[18]), .IN4(n13), .IN5(n87), .Q(
        n35) );
  AO22X1 U86 ( .IN1(A[15]), .IN2(n10), .IN3(A[16]), .IN4(n9), .Q(n87) );
  AO221X1 U87 ( .IN1(A[13]), .IN2(n12), .IN3(A[14]), .IN4(n13), .IN5(n88), .Q(
        n29) );
  AO22X1 U88 ( .IN1(A[11]), .IN2(n10), .IN3(A[12]), .IN4(n9), .Q(n88) );
  AO221X1 U89 ( .IN1(n12), .IN2(A[21]), .IN3(n13), .IN4(A[22]), .IN5(n89), .Q(
        n32) );
  AO22X1 U90 ( .IN1(n10), .IN2(A[19]), .IN3(A[20]), .IN4(n9), .Q(n89) );
  AO222X1 U91 ( .IN1(n21), .IN2(n82), .IN3(n19), .IN4(n37), .IN5(n23), .IN6(
        n39), .Q(B[10]) );
  AO221X1 U92 ( .IN1(A[16]), .IN2(n12), .IN3(A[17]), .IN4(n13), .IN5(n90), .Q(
        n39) );
  AO22X1 U93 ( .IN1(A[14]), .IN2(n10), .IN3(A[15]), .IN4(n9), .Q(n90) );
  NOR2X0 U94 ( .IN1(n91), .IN2(n81), .QN(n23) );
  AO221X1 U95 ( .IN1(A[12]), .IN2(n12), .IN3(A[13]), .IN4(n13), .IN5(n92), .Q(
        n37) );
  AO22X1 U96 ( .IN1(A[10]), .IN2(n10), .IN3(A[11]), .IN4(n9), .Q(n92) );
  NOR2X0 U97 ( .IN1(n54), .IN2(SH[7]), .QN(n19) );
  AO21X1 U98 ( .IN1(A[22]), .IN2(n11), .IN3(n9), .Q(n84) );
  AO221X1 U99 ( .IN1(A[20]), .IN2(n12), .IN3(n13), .IN4(A[21]), .IN5(n93), .Q(
        n40) );
  AO22X1 U100 ( .IN1(n10), .IN2(A[18]), .IN3(A[19]), .IN4(n9), .Q(n93) );
  NOR2X0 U101 ( .IN1(n81), .IN2(n65), .QN(n21) );
  NAND2X0 U102 ( .IN1(n66), .IN2(n1), .QN(n81) );
  NOR2X0 U103 ( .IN1(SH[7]), .IN2(n94), .QN(B[0]) );
  OA21X1 U104 ( .IN1(n95), .IN2(n54), .IN3(n96), .Q(n94) );
  MUX21X1 U105 ( .IN1(n83), .IN2(n97), .S(n66), .Q(n96) );
  AOI222X1 U106 ( .IN1(n46), .IN2(n3), .IN3(n25), .IN4(n58), .IN5(n27), .IN6(
        n59), .QN(n97) );
  NOR2X0 U107 ( .IN1(n8), .IN2(n65), .QN(n59) );
  AO221X1 U108 ( .IN1(A[14]), .IN2(n12), .IN3(A[15]), .IN4(n13), .IN5(n98), 
        .Q(n27) );
  AO22X1 U109 ( .IN1(A[12]), .IN2(n10), .IN3(A[13]), .IN4(n9), .Q(n98) );
  NOR2X0 U110 ( .IN1(n65), .IN2(SH[2]), .QN(n58) );
  AO221X1 U111 ( .IN1(A[10]), .IN2(n12), .IN3(A[11]), .IN4(n13), .IN5(n99), 
        .Q(n25) );
  AO22X1 U112 ( .IN1(A[8]), .IN2(n10), .IN3(A[9]), .IN4(n9), .Q(n99) );
  NAND2X0 U113 ( .IN1(n65), .IN2(SH[2]), .QN(n91) );
  AO221X1 U114 ( .IN1(A[6]), .IN2(n12), .IN3(A[7]), .IN4(n13), .IN5(n100), .Q(
        n46) );
  AO22X1 U115 ( .IN1(A[4]), .IN2(n10), .IN3(A[5]), .IN4(n9), .Q(n100) );
  NAND2X0 U116 ( .IN1(n65), .IN2(n26), .QN(n83) );
  MUX21X1 U117 ( .IN1(n49), .IN2(n48), .S(n8), .Q(n26) );
  AO221X1 U118 ( .IN1(A[18]), .IN2(n12), .IN3(n13), .IN4(A[19]), .IN5(n101), 
        .Q(n48) );
  AO22X1 U119 ( .IN1(A[16]), .IN2(n10), .IN3(A[17]), .IN4(n9), .Q(n101) );
  AO21X1 U120 ( .IN1(n10), .IN2(A[20]), .IN3(n13), .Q(n102) );
  NAND3X0 U121 ( .IN1(n66), .IN2(n8), .IN3(n65), .QN(n54) );
  NOR2X0 U122 ( .IN1(SH[3]), .IN2(n103), .QN(n65) );
  NOR2X0 U123 ( .IN1(SH[4]), .IN2(n103), .QN(n66) );
  OR2X1 U124 ( .IN1(SH[5]), .IN2(SH[6]), .Q(n103) );
  OA221X1 U125 ( .IN1(n79), .IN2(n16), .IN3(n78), .IN4(n17), .IN5(n104), .Q(
        n95) );
  AOI22X1 U126 ( .IN1(A[1]), .IN2(n9), .IN3(A[0]), .IN4(n10), .QN(n104) );
  NAND2X0 U127 ( .IN1(n14), .IN2(n11), .QN(n55) );
  NAND2X0 U128 ( .IN1(SH[0]), .IN2(n11), .QN(n56) );
  NAND2X0 U129 ( .IN1(SH[1]), .IN2(n14), .QN(n78) );
  NAND2X0 U130 ( .IN1(SH[0]), .IN2(SH[1]), .QN(n79) );
endmodule


module booth_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND3X0 U3 ( .IN1(n65), .IN2(n66), .IN3(n1), .QN(n69) );
  AO221X1 U4 ( .IN1(A[21]), .IN2(SH[0]), .IN3(A[22]), .IN4(SH[1]), .IN5(n102), 
        .Q(n49) );
  INVX0 U5 ( .INP(n55), .ZN(n10) );
  INVX0 U6 ( .INP(n68), .ZN(n7) );
  INVX0 U7 ( .INP(n75), .ZN(n4) );
  INVX0 U8 ( .INP(n80), .ZN(n5) );
  INVX0 U9 ( .INP(n82), .ZN(n6) );
  INVX0 U10 ( .INP(n91), .ZN(n3) );
  INVX0 U11 ( .INP(n56), .ZN(n9) );
  INVX0 U12 ( .INP(n78), .ZN(n12) );
  AND2X1 U13 ( .IN1(n21), .IN2(SH[2]), .Q(n31) );
  MUX21X1 U14 ( .IN1(n40), .IN2(n84), .S(SH[2]), .Q(n82) );
  MUX21X1 U15 ( .IN1(n32), .IN2(n10), .S(SH[2]), .Q(n80) );
  INVX0 U16 ( .INP(n79), .ZN(n13) );
  INVX0 U17 ( .INP(n66), .ZN(n2) );
  INVX0 U18 ( .INP(SH[7]), .ZN(n1) );
  INVX0 U19 ( .INP(SH[0]), .ZN(n14) );
  INVX0 U20 ( .INP(SH[1]), .ZN(n11) );
  INVX0 U21 ( .INP(A[1]), .ZN(n18) );
  INVX0 U22 ( .INP(A[4]), .ZN(n15) );
  INVX0 U23 ( .INP(A[3]), .ZN(n16) );
  INVX0 U24 ( .INP(A[2]), .ZN(n17) );
  INVX0 U25 ( .INP(SH[2]), .ZN(n8) );
  AO222X1 U26 ( .IN1(n19), .IN2(n20), .IN3(n21), .IN4(n22), .IN5(n23), .IN6(
        n24), .Q(B[9]) );
  AO222X1 U27 ( .IN1(n19), .IN2(n25), .IN3(n21), .IN4(n26), .IN5(n23), .IN6(
        n27), .Q(B[8]) );
  AO221X1 U28 ( .IN1(n19), .IN2(n28), .IN3(n23), .IN4(n29), .IN5(n30), .Q(B[7]) );
  AO222X1 U29 ( .IN1(n31), .IN2(n32), .IN3(n33), .IN4(n10), .IN5(n34), .IN6(
        n35), .Q(n30) );
  AO221X1 U30 ( .IN1(n19), .IN2(n36), .IN3(n23), .IN4(n37), .IN5(n38), .Q(B[6]) );
  AO222X1 U31 ( .IN1(n34), .IN2(n39), .IN3(n31), .IN4(n40), .IN5(n7), .IN6(n41), .Q(n38) );
  AO221X1 U32 ( .IN1(n19), .IN2(n42), .IN3(n23), .IN4(n20), .IN5(n43), .Q(B[5]) );
  AO222X1 U33 ( .IN1(n31), .IN2(n44), .IN3(n33), .IN4(n45), .IN5(n34), .IN6(
        n24), .Q(n43) );
  AO221X1 U34 ( .IN1(n19), .IN2(n46), .IN3(n23), .IN4(n25), .IN5(n47), .Q(B[4]) );
  AO222X1 U35 ( .IN1(n31), .IN2(n48), .IN3(n33), .IN4(n49), .IN5(n34), .IN6(
        n27), .Q(n47) );
  AND2X1 U36 ( .IN1(n41), .IN2(n8), .Q(n33) );
  NOR2X0 U37 ( .IN1(n50), .IN2(SH[7]), .QN(n41) );
  NOR2X0 U38 ( .IN1(SH[7]), .IN2(n51), .QN(B[3]) );
  OA222X1 U39 ( .IN1(n52), .IN2(n2), .IN3(n5), .IN4(n50), .IN5(n53), .IN6(n54), 
        .Q(n51) );
  OA221X1 U40 ( .IN1(n55), .IN2(n16), .IN3(n56), .IN4(n15), .IN5(n57), .Q(n53)
         );
  AOI22X1 U41 ( .IN1(n12), .IN2(A[5]), .IN3(n13), .IN4(A[6]), .QN(n57) );
  AOI222X1 U42 ( .IN1(n28), .IN2(n3), .IN3(n29), .IN4(n58), .IN5(n35), .IN6(
        n59), .QN(n52) );
  AO221X1 U43 ( .IN1(A[9]), .IN2(n12), .IN3(A[10]), .IN4(n13), .IN5(n60), .Q(
        n28) );
  AO22X1 U44 ( .IN1(A[7]), .IN2(n10), .IN3(A[8]), .IN4(n9), .Q(n60) );
  NOR2X0 U45 ( .IN1(SH[7]), .IN2(n61), .QN(B[2]) );
  OA222X1 U46 ( .IN1(n62), .IN2(n2), .IN3(n6), .IN4(n50), .IN5(n63), .IN6(n54), 
        .Q(n61) );
  OA221X1 U47 ( .IN1(n55), .IN2(n17), .IN3(n56), .IN4(n16), .IN5(n64), .Q(n63)
         );
  AOI22X1 U48 ( .IN1(n12), .IN2(A[4]), .IN3(n13), .IN4(A[5]), .QN(n64) );
  NAND2X0 U49 ( .IN1(n65), .IN2(n2), .QN(n50) );
  AOI222X1 U50 ( .IN1(n36), .IN2(n3), .IN3(n37), .IN4(n58), .IN5(n39), .IN6(
        n59), .QN(n62) );
  AO221X1 U51 ( .IN1(A[8]), .IN2(n12), .IN3(A[9]), .IN4(n13), .IN5(n67), .Q(
        n36) );
  AO22X1 U52 ( .IN1(A[6]), .IN2(n10), .IN3(A[7]), .IN4(n9), .Q(n67) );
  AND2X1 U53 ( .IN1(n10), .IN2(n19), .Q(B[23]) );
  NOR2X0 U54 ( .IN1(n68), .IN2(n69), .QN(B[22]) );
  AND2X1 U55 ( .IN1(n45), .IN2(n19), .Q(B[21]) );
  AND2X1 U56 ( .IN1(n49), .IN2(n19), .Q(B[20]) );
  OA21X1 U57 ( .IN1(n70), .IN2(n71), .IN3(n1), .Q(B[1]) );
  MUX21X1 U58 ( .IN1(n4), .IN2(n72), .S(n66), .Q(n71) );
  AO222X1 U59 ( .IN1(n59), .IN2(n24), .IN3(n58), .IN4(n20), .IN5(n3), .IN6(n42), .Q(n72) );
  AO221X1 U60 ( .IN1(A[7]), .IN2(n12), .IN3(A[8]), .IN4(n13), .IN5(n73), .Q(
        n42) );
  AO22X1 U61 ( .IN1(A[5]), .IN2(n10), .IN3(A[6]), .IN4(n9), .Q(n73) );
  AO221X1 U62 ( .IN1(A[11]), .IN2(n12), .IN3(A[12]), .IN4(n13), .IN5(n74), .Q(
        n20) );
  AO22X1 U63 ( .IN1(A[9]), .IN2(n10), .IN3(A[10]), .IN4(n9), .Q(n74) );
  NOR2X0 U64 ( .IN1(n76), .IN2(n54), .QN(n70) );
  OA221X1 U65 ( .IN1(n55), .IN2(n18), .IN3(n56), .IN4(n17), .IN5(n77), .Q(n76)
         );
  OA22X1 U66 ( .IN1(n78), .IN2(n16), .IN3(n79), .IN4(n15), .Q(n77) );
  NOR2X0 U67 ( .IN1(n5), .IN2(n69), .QN(B[19]) );
  NOR2X0 U68 ( .IN1(n6), .IN2(n69), .QN(B[18]) );
  NOR2X0 U69 ( .IN1(n81), .IN2(n75), .QN(B[17]) );
  NAND2X0 U70 ( .IN1(n65), .IN2(n22), .QN(n75) );
  MUX21X1 U71 ( .IN1(n45), .IN2(n44), .S(n8), .Q(n22) );
  NOR2X0 U72 ( .IN1(n81), .IN2(n83), .QN(B[16]) );
  AO222X1 U73 ( .IN1(n19), .IN2(n35), .IN3(n34), .IN4(n10), .IN5(n23), .IN6(
        n32), .Q(B[15]) );
  AO222X1 U74 ( .IN1(n7), .IN2(n21), .IN3(n19), .IN4(n39), .IN5(n23), .IN6(n40), .Q(B[14]) );
  NAND2X0 U75 ( .IN1(n84), .IN2(n8), .QN(n68) );
  AO222X1 U76 ( .IN1(n19), .IN2(n24), .IN3(n34), .IN4(n45), .IN5(n23), .IN6(
        n44), .Q(B[13]) );
  AO221X1 U77 ( .IN1(A[19]), .IN2(n12), .IN3(A[20]), .IN4(n13), .IN5(n85), .Q(
        n44) );
  AO22X1 U78 ( .IN1(A[17]), .IN2(n10), .IN3(A[18]), .IN4(n9), .Q(n85) );
  AO221X1 U79 ( .IN1(A[22]), .IN2(n9), .IN3(A[21]), .IN4(n14), .IN5(n12), .Q(
        n45) );
  AO221X1 U80 ( .IN1(A[15]), .IN2(n12), .IN3(A[16]), .IN4(n13), .IN5(n86), .Q(
        n24) );
  AO22X1 U81 ( .IN1(A[13]), .IN2(n10), .IN3(A[14]), .IN4(n9), .Q(n86) );
  AO222X1 U82 ( .IN1(n19), .IN2(n27), .IN3(n34), .IN4(n49), .IN5(n23), .IN6(
        n48), .Q(B[12]) );
  AND2X1 U83 ( .IN1(n21), .IN2(n8), .Q(n34) );
  AO222X1 U84 ( .IN1(n21), .IN2(n80), .IN3(n19), .IN4(n29), .IN5(n23), .IN6(
        n35), .Q(B[11]) );
  AO221X1 U85 ( .IN1(A[17]), .IN2(n12), .IN3(A[18]), .IN4(n13), .IN5(n87), .Q(
        n35) );
  AO22X1 U86 ( .IN1(A[15]), .IN2(n10), .IN3(A[16]), .IN4(n9), .Q(n87) );
  AO221X1 U87 ( .IN1(A[13]), .IN2(n12), .IN3(A[14]), .IN4(n13), .IN5(n88), .Q(
        n29) );
  AO22X1 U88 ( .IN1(A[11]), .IN2(n10), .IN3(A[12]), .IN4(n9), .Q(n88) );
  AO221X1 U89 ( .IN1(n12), .IN2(A[21]), .IN3(n13), .IN4(A[22]), .IN5(n89), .Q(
        n32) );
  AO22X1 U90 ( .IN1(n10), .IN2(A[19]), .IN3(A[20]), .IN4(n9), .Q(n89) );
  AO222X1 U91 ( .IN1(n21), .IN2(n82), .IN3(n19), .IN4(n37), .IN5(n23), .IN6(
        n39), .Q(B[10]) );
  AO221X1 U92 ( .IN1(A[16]), .IN2(n12), .IN3(A[17]), .IN4(n13), .IN5(n90), .Q(
        n39) );
  AO22X1 U93 ( .IN1(A[14]), .IN2(n10), .IN3(A[15]), .IN4(n9), .Q(n90) );
  NOR2X0 U94 ( .IN1(n91), .IN2(n81), .QN(n23) );
  AO221X1 U95 ( .IN1(A[12]), .IN2(n12), .IN3(A[13]), .IN4(n13), .IN5(n92), .Q(
        n37) );
  AO22X1 U96 ( .IN1(A[10]), .IN2(n10), .IN3(A[11]), .IN4(n9), .Q(n92) );
  NOR2X0 U97 ( .IN1(n54), .IN2(SH[7]), .QN(n19) );
  AO21X1 U98 ( .IN1(A[22]), .IN2(n11), .IN3(n9), .Q(n84) );
  AO221X1 U99 ( .IN1(A[20]), .IN2(n12), .IN3(n13), .IN4(A[21]), .IN5(n93), .Q(
        n40) );
  AO22X1 U100 ( .IN1(n10), .IN2(A[18]), .IN3(A[19]), .IN4(n9), .Q(n93) );
  NOR2X0 U101 ( .IN1(n81), .IN2(n65), .QN(n21) );
  NAND2X0 U102 ( .IN1(n66), .IN2(n1), .QN(n81) );
  NOR2X0 U103 ( .IN1(SH[7]), .IN2(n94), .QN(B[0]) );
  OA21X1 U104 ( .IN1(n95), .IN2(n54), .IN3(n96), .Q(n94) );
  MUX21X1 U105 ( .IN1(n83), .IN2(n97), .S(n66), .Q(n96) );
  AOI222X1 U106 ( .IN1(n46), .IN2(n3), .IN3(n25), .IN4(n58), .IN5(n27), .IN6(
        n59), .QN(n97) );
  NOR2X0 U107 ( .IN1(n8), .IN2(n65), .QN(n59) );
  AO221X1 U108 ( .IN1(A[14]), .IN2(n12), .IN3(A[15]), .IN4(n13), .IN5(n98), 
        .Q(n27) );
  AO22X1 U109 ( .IN1(A[12]), .IN2(n10), .IN3(A[13]), .IN4(n9), .Q(n98) );
  NOR2X0 U110 ( .IN1(n65), .IN2(SH[2]), .QN(n58) );
  AO221X1 U111 ( .IN1(A[10]), .IN2(n12), .IN3(A[11]), .IN4(n13), .IN5(n99), 
        .Q(n25) );
  AO22X1 U112 ( .IN1(A[8]), .IN2(n10), .IN3(A[9]), .IN4(n9), .Q(n99) );
  NAND2X0 U113 ( .IN1(n65), .IN2(SH[2]), .QN(n91) );
  AO221X1 U114 ( .IN1(A[6]), .IN2(n12), .IN3(A[7]), .IN4(n13), .IN5(n100), .Q(
        n46) );
  AO22X1 U115 ( .IN1(A[4]), .IN2(n10), .IN3(A[5]), .IN4(n9), .Q(n100) );
  NAND2X0 U116 ( .IN1(n65), .IN2(n26), .QN(n83) );
  MUX21X1 U117 ( .IN1(n49), .IN2(n48), .S(n8), .Q(n26) );
  AO221X1 U118 ( .IN1(A[18]), .IN2(n12), .IN3(n13), .IN4(A[19]), .IN5(n101), 
        .Q(n48) );
  AO22X1 U119 ( .IN1(A[16]), .IN2(n10), .IN3(A[17]), .IN4(n9), .Q(n101) );
  AO21X1 U120 ( .IN1(n10), .IN2(A[20]), .IN3(n13), .Q(n102) );
  NAND3X0 U121 ( .IN1(n66), .IN2(n8), .IN3(n65), .QN(n54) );
  NOR2X0 U122 ( .IN1(SH[3]), .IN2(n103), .QN(n65) );
  NOR2X0 U123 ( .IN1(SH[4]), .IN2(n103), .QN(n66) );
  OR2X1 U124 ( .IN1(SH[5]), .IN2(SH[6]), .Q(n103) );
  OA221X1 U125 ( .IN1(n79), .IN2(n16), .IN3(n78), .IN4(n17), .IN5(n104), .Q(
        n95) );
  AOI22X1 U126 ( .IN1(A[1]), .IN2(n9), .IN3(A[0]), .IN4(n10), .QN(n104) );
  NAND2X0 U127 ( .IN1(n14), .IN2(n11), .QN(n55) );
  NAND2X0 U128 ( .IN1(SH[0]), .IN2(n11), .QN(n56) );
  NAND2X0 U129 ( .IN1(SH[1]), .IN2(n14), .QN(n78) );
  NAND2X0 U130 ( .IN1(SH[0]), .IN2(SH[1]), .QN(n79) );
endmodule


module booth ( clk, reset, combined_a, combined_b, combined_negative_b, 
        product_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_exponent_a, add_difference, 
        add_zero_flag, add_greater_flag, add_lesser_flag, add_fraction_a, 
        add_fraction_b, add_combined_a_o, add_combined_b_o, new_add_exponent_o, 
        add_sign_a2, add_sign_b2, add_sign_a3, add_sign_b3, s, s2, 
        add_greater_flag2 );
  input [24:0] combined_a;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [7:0] add_exponent_a;
  input [7:0] add_difference;
  input [22:0] add_fraction_a;
  input [22:0] add_fraction_b;
  output [23:0] add_combined_a_o;
  output [23:0] add_combined_b_o;
  output [7:0] new_add_exponent_o;
  input clk, reset, new_sign, add_zero_flag, add_greater_flag, add_lesser_flag,
         add_sign_a2, add_sign_b2, s;
  output new_sign2, add_sign_a3, add_sign_b3, s2, add_greater_flag2;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, n15, n16,
         n17, n18, n19, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;
  wire   [50:0] product;
  wire   [7:0] new_add_exponent;
  wire   [23:0] add_combined_a;
  wire   [23:0] add_combined_b;
  assign product_o[25] = 1'b0;
  assign N12 = combined_a[1];
  assign N13 = combined_a[2];
  assign N14 = combined_a[3];
  assign N15 = combined_a[4];
  assign N16 = combined_a[5];
  assign N17 = combined_a[6];
  assign N18 = combined_a[7];
  assign N19 = combined_a[8];
  assign N20 = combined_a[9];
  assign N21 = combined_a[10];
  assign N22 = combined_a[11];
  assign N23 = combined_a[12];
  assign N24 = combined_a[13];
  assign N25 = combined_a[14];
  assign N26 = combined_a[15];
  assign N27 = combined_a[16];
  assign N28 = combined_a[17];
  assign N29 = combined_a[18];
  assign N30 = combined_a[19];
  assign N31 = combined_a[20];
  assign N32 = combined_a[21];
  assign N33 = combined_a[22];
  assign N34 = combined_a[23];
  assign N36 = combined_negative_b[0];
  assign N37 = combined_negative_b[1];
  assign N38 = combined_negative_b[2];
  assign N39 = combined_negative_b[3];
  assign N40 = combined_negative_b[4];
  assign N41 = combined_negative_b[5];
  assign N42 = combined_negative_b[6];
  assign N43 = combined_negative_b[7];
  assign N44 = combined_negative_b[8];
  assign N45 = combined_negative_b[9];
  assign N46 = combined_negative_b[10];
  assign N47 = combined_negative_b[11];
  assign N48 = combined_negative_b[12];
  assign N49 = combined_negative_b[13];
  assign N50 = combined_negative_b[14];
  assign N51 = combined_negative_b[15];
  assign N52 = combined_negative_b[16];
  assign N53 = combined_negative_b[17];
  assign N54 = combined_negative_b[18];
  assign N55 = combined_negative_b[19];
  assign N56 = combined_negative_b[20];
  assign N57 = combined_negative_b[21];
  assign N58 = combined_negative_b[22];
  assign N59 = combined_negative_b[23];
  assign N60 = combined_negative_b[24];

  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n35), .Q(new_sign2)
         );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n35), .Q(s2) );
  DFFARX1 \product_o_reg[50]  ( .D(product[50]), .CLK(clk), .RSTB(n34), .Q(
        product_o[50]) );
  DFFARX1 \product_o_reg[49]  ( .D(product[49]), .CLK(clk), .RSTB(n34), .Q(
        product_o[49]) );
  DFFARX1 \product_o_reg[48]  ( .D(product[48]), .CLK(clk), .RSTB(n34), .Q(
        product_o[48]) );
  DFFARX1 \product_o_reg[47]  ( .D(product[47]), .CLK(clk), .RSTB(n34), .Q(
        product_o[47]) );
  DFFARX1 \product_o_reg[46]  ( .D(product[46]), .CLK(clk), .RSTB(n34), .Q(
        product_o[46]) );
  DFFARX1 \product_o_reg[45]  ( .D(product[45]), .CLK(clk), .RSTB(n34), .Q(
        product_o[45]) );
  DFFARX1 \product_o_reg[44]  ( .D(product[44]), .CLK(clk), .RSTB(n34), .Q(
        product_o[44]) );
  DFFARX1 \product_o_reg[43]  ( .D(product[43]), .CLK(clk), .RSTB(n34), .Q(
        product_o[43]) );
  DFFARX1 \product_o_reg[42]  ( .D(product[42]), .CLK(clk), .RSTB(n34), .Q(
        product_o[42]) );
  DFFARX1 \product_o_reg[41]  ( .D(product[41]), .CLK(clk), .RSTB(n34), .Q(
        product_o[41]) );
  DFFARX1 \product_o_reg[40]  ( .D(product[40]), .CLK(clk), .RSTB(n34), .Q(
        product_o[40]) );
  DFFARX1 \product_o_reg[39]  ( .D(product[39]), .CLK(clk), .RSTB(n34), .Q(
        product_o[39]) );
  DFFARX1 \product_o_reg[38]  ( .D(product[38]), .CLK(clk), .RSTB(n33), .Q(
        product_o[38]) );
  DFFARX1 \product_o_reg[37]  ( .D(product[37]), .CLK(clk), .RSTB(n33), .Q(
        product_o[37]) );
  DFFARX1 \product_o_reg[36]  ( .D(product[36]), .CLK(clk), .RSTB(n33), .Q(
        product_o[36]) );
  DFFARX1 \product_o_reg[35]  ( .D(product[35]), .CLK(clk), .RSTB(n33), .Q(
        product_o[35]) );
  DFFARX1 \product_o_reg[34]  ( .D(product[34]), .CLK(clk), .RSTB(n33), .Q(
        product_o[34]) );
  DFFARX1 \product_o_reg[33]  ( .D(product[33]), .CLK(clk), .RSTB(n33), .Q(
        product_o[33]) );
  DFFARX1 \product_o_reg[32]  ( .D(product[32]), .CLK(clk), .RSTB(n33), .Q(
        product_o[32]) );
  DFFARX1 \product_o_reg[31]  ( .D(product[31]), .CLK(clk), .RSTB(n33), .Q(
        product_o[31]) );
  DFFARX1 \product_o_reg[30]  ( .D(product[30]), .CLK(clk), .RSTB(n33), .Q(
        product_o[30]) );
  DFFARX1 \product_o_reg[29]  ( .D(product[29]), .CLK(clk), .RSTB(n33), .Q(
        product_o[29]) );
  DFFARX1 \product_o_reg[28]  ( .D(product[28]), .CLK(clk), .RSTB(n33), .Q(
        product_o[28]) );
  DFFARX1 \product_o_reg[27]  ( .D(product[27]), .CLK(clk), .RSTB(n33), .Q(
        product_o[27]) );
  DFFARX1 \product_o_reg[26]  ( .D(product[26]), .CLK(clk), .RSTB(n32), .Q(
        product_o[26]) );
  DFFARX1 \product_o_reg[24]  ( .D(product[24]), .CLK(clk), .RSTB(n32), .Q(
        product_o[24]) );
  DFFARX1 \product_o_reg[23]  ( .D(product[23]), .CLK(clk), .RSTB(n32), .Q(
        product_o[23]) );
  DFFARX1 \product_o_reg[22]  ( .D(product[22]), .CLK(clk), .RSTB(n32), .Q(
        product_o[22]) );
  DFFARX1 \product_o_reg[21]  ( .D(product[21]), .CLK(clk), .RSTB(n32), .Q(
        product_o[21]) );
  DFFARX1 \product_o_reg[20]  ( .D(product[20]), .CLK(clk), .RSTB(n32), .Q(
        product_o[20]) );
  DFFARX1 \product_o_reg[19]  ( .D(product[19]), .CLK(clk), .RSTB(n32), .Q(
        product_o[19]) );
  DFFARX1 \product_o_reg[18]  ( .D(product[18]), .CLK(clk), .RSTB(n32), .Q(
        product_o[18]) );
  DFFARX1 \product_o_reg[17]  ( .D(product[17]), .CLK(clk), .RSTB(n32), .Q(
        product_o[17]) );
  DFFARX1 \product_o_reg[16]  ( .D(product[16]), .CLK(clk), .RSTB(n32), .Q(
        product_o[16]) );
  DFFARX1 \product_o_reg[15]  ( .D(product[15]), .CLK(clk), .RSTB(n32), .Q(
        product_o[15]) );
  DFFARX1 \product_o_reg[14]  ( .D(product[14]), .CLK(clk), .RSTB(n31), .Q(
        product_o[14]) );
  DFFARX1 \product_o_reg[13]  ( .D(product[13]), .CLK(clk), .RSTB(n31), .Q(
        product_o[13]) );
  DFFARX1 \product_o_reg[12]  ( .D(product[12]), .CLK(clk), .RSTB(n31), .Q(
        product_o[12]) );
  DFFARX1 \product_o_reg[11]  ( .D(product[11]), .CLK(clk), .RSTB(n31), .Q(
        product_o[11]) );
  DFFARX1 \product_o_reg[10]  ( .D(product[10]), .CLK(clk), .RSTB(n31), .Q(
        product_o[10]) );
  DFFARX1 \product_o_reg[9]  ( .D(product[9]), .CLK(clk), .RSTB(n31), .Q(
        product_o[9]) );
  DFFARX1 \product_o_reg[8]  ( .D(product[8]), .CLK(clk), .RSTB(n31), .Q(
        product_o[8]) );
  DFFARX1 \product_o_reg[7]  ( .D(product[7]), .CLK(clk), .RSTB(n31), .Q(
        product_o[7]) );
  DFFARX1 \product_o_reg[6]  ( .D(product[6]), .CLK(clk), .RSTB(n31), .Q(
        product_o[6]) );
  DFFARX1 \product_o_reg[5]  ( .D(product[5]), .CLK(clk), .RSTB(n31), .Q(
        product_o[5]) );
  DFFARX1 \product_o_reg[4]  ( .D(product[4]), .CLK(clk), .RSTB(n31), .Q(
        product_o[4]) );
  DFFARX1 \product_o_reg[3]  ( .D(product[3]), .CLK(clk), .RSTB(n31), .Q(
        product_o[3]) );
  DFFARX1 \product_o_reg[2]  ( .D(product[2]), .CLK(clk), .RSTB(n30), .Q(
        product_o[2]) );
  DFFARX1 \product_o_reg[1]  ( .D(n13), .CLK(clk), .RSTB(n30), .Q(product_o[1]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n30), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n22), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n22), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n22), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n22), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n22), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n22), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n22), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(combined_b[7]), .CLK(clk), .RSTB(n22), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(combined_b[6]), .CLK(clk), .RSTB(n22), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(combined_b[5]), .CLK(clk), .RSTB(n22), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(combined_b[4]), .CLK(clk), .RSTB(n35), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(combined_b[3]), .CLK(clk), .RSTB(n35), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(combined_b[2]), .CLK(clk), .RSTB(n29), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n29), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n29), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(N60), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(N59), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(N58), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(N57), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(N56), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(N55), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(N54), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(N53), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(N52), .CLK(clk), .RSTB(n29), .Q(
        combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(N51), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(N50), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(N49), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(N48), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(N47), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(N46), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(N45), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(N44), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(N43), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(N42), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(N41), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(N40), .CLK(clk), .RSTB(n28), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(N39), .CLK(clk), .RSTB(n27), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(N38), .CLK(clk), .RSTB(n27), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(N37), .CLK(clk), .RSTB(n27), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(N36), .CLK(clk), .RSTB(n27), .Q(
        combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n27), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n26), 
        .Q(new_exponent2[0]) );
  DFFARX1 add_sign_b3_reg ( .D(add_sign_b2), .CLK(clk), .RSTB(n26), .Q(
        add_sign_b3) );
  DFFARX1 add_greater_flag2_reg ( .D(add_greater_flag), .CLK(clk), .RSTB(n26), 
        .Q(add_greater_flag2) );
  DFFARX1 \new_add_exponent_o_reg[7]  ( .D(new_add_exponent[7]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[7]) );
  DFFARX1 \new_add_exponent_o_reg[6]  ( .D(new_add_exponent[6]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[6]) );
  DFFARX1 \new_add_exponent_o_reg[5]  ( .D(new_add_exponent[5]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[5]) );
  DFFARX1 \new_add_exponent_o_reg[4]  ( .D(new_add_exponent[4]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[4]) );
  DFFARX1 \new_add_exponent_o_reg[3]  ( .D(new_add_exponent[3]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[3]) );
  DFFARX1 \new_add_exponent_o_reg[2]  ( .D(new_add_exponent[2]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[2]) );
  DFFARX1 \new_add_exponent_o_reg[1]  ( .D(new_add_exponent[1]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[1]) );
  DFFARX1 \new_add_exponent_o_reg[0]  ( .D(new_add_exponent[0]), .CLK(clk), 
        .RSTB(n26), .Q(new_add_exponent_o[0]) );
  DFFARX1 \add_combined_a_o_reg[23]  ( .D(add_combined_a[23]), .CLK(clk), 
        .RSTB(n26), .Q(add_combined_a_o[23]) );
  DFFARX1 \add_combined_a_o_reg[22]  ( .D(add_combined_a[22]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[22]) );
  DFFARX1 \add_combined_a_o_reg[21]  ( .D(add_combined_a[21]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[21]) );
  DFFARX1 \add_combined_a_o_reg[20]  ( .D(add_combined_a[20]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[20]) );
  DFFARX1 \add_combined_a_o_reg[19]  ( .D(add_combined_a[19]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[19]) );
  DFFARX1 \add_combined_a_o_reg[18]  ( .D(add_combined_a[18]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[18]) );
  DFFARX1 \add_combined_a_o_reg[17]  ( .D(add_combined_a[17]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[17]) );
  DFFARX1 \add_combined_a_o_reg[16]  ( .D(add_combined_a[16]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[16]) );
  DFFARX1 \add_combined_a_o_reg[15]  ( .D(add_combined_a[15]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[15]) );
  DFFARX1 \add_combined_a_o_reg[14]  ( .D(add_combined_a[14]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[14]) );
  DFFARX1 \add_combined_a_o_reg[13]  ( .D(add_combined_a[13]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[13]) );
  DFFARX1 \add_combined_a_o_reg[12]  ( .D(add_combined_a[12]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[12]) );
  DFFARX1 \add_combined_a_o_reg[11]  ( .D(add_combined_a[11]), .CLK(clk), 
        .RSTB(n25), .Q(add_combined_a_o[11]) );
  DFFARX1 \add_combined_a_o_reg[10]  ( .D(add_combined_a[10]), .CLK(clk), 
        .RSTB(n24), .Q(add_combined_a_o[10]) );
  DFFARX1 \add_combined_a_o_reg[9]  ( .D(add_combined_a[9]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[9]) );
  DFFARX1 \add_combined_a_o_reg[8]  ( .D(add_combined_a[8]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[8]) );
  DFFARX1 \add_combined_a_o_reg[7]  ( .D(add_combined_a[7]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[7]) );
  DFFARX1 \add_combined_a_o_reg[6]  ( .D(add_combined_a[6]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[6]) );
  DFFARX1 \add_combined_a_o_reg[5]  ( .D(add_combined_a[5]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[5]) );
  DFFARX1 \add_combined_a_o_reg[4]  ( .D(add_combined_a[4]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[4]) );
  DFFARX1 \add_combined_a_o_reg[3]  ( .D(add_combined_a[3]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[3]) );
  DFFARX1 \add_combined_a_o_reg[2]  ( .D(add_combined_a[2]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[2]) );
  DFFARX1 \add_combined_a_o_reg[1]  ( .D(add_combined_a[1]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[1]) );
  DFFARX1 \add_combined_a_o_reg[0]  ( .D(add_combined_a[0]), .CLK(clk), .RSTB(
        n24), .Q(add_combined_a_o[0]) );
  DFFARX1 \add_combined_b_o_reg[23]  ( .D(add_combined_b[23]), .CLK(clk), 
        .RSTB(n24), .Q(add_combined_b_o[23]) );
  DFFARX1 \add_combined_b_o_reg[22]  ( .D(add_combined_b[22]), .CLK(clk), 
        .RSTB(n21), .Q(add_combined_b_o[22]) );
  DFFARX1 \add_combined_b_o_reg[21]  ( .D(add_combined_b[21]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[21]) );
  DFFARX1 \add_combined_b_o_reg[20]  ( .D(add_combined_b[20]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[20]) );
  DFFARX1 \add_combined_b_o_reg[19]  ( .D(add_combined_b[19]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[19]) );
  DFFARX1 \add_combined_b_o_reg[18]  ( .D(add_combined_b[18]), .CLK(clk), 
        .RSTB(n21), .Q(add_combined_b_o[18]) );
  DFFARX1 \add_combined_b_o_reg[17]  ( .D(add_combined_b[17]), .CLK(clk), 
        .RSTB(n21), .Q(add_combined_b_o[17]) );
  DFFARX1 \add_combined_b_o_reg[16]  ( .D(add_combined_b[16]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[16]) );
  DFFARX1 \add_combined_b_o_reg[15]  ( .D(add_combined_b[15]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[15]) );
  DFFARX1 \add_combined_b_o_reg[14]  ( .D(add_combined_b[14]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[14]) );
  DFFARX1 \add_combined_b_o_reg[13]  ( .D(add_combined_b[13]), .CLK(clk), 
        .RSTB(n30), .Q(add_combined_b_o[13]) );
  DFFARX1 \add_combined_b_o_reg[12]  ( .D(add_combined_b[12]), .CLK(clk), 
        .RSTB(n32), .Q(add_combined_b_o[12]) );
  DFFARX1 \add_combined_b_o_reg[11]  ( .D(add_combined_b[11]), .CLK(clk), 
        .RSTB(n35), .Q(add_combined_b_o[11]) );
  DFFARX1 \add_combined_b_o_reg[10]  ( .D(add_combined_b[10]), .CLK(clk), 
        .RSTB(n23), .Q(add_combined_b_o[10]) );
  DFFARX1 \add_combined_b_o_reg[9]  ( .D(add_combined_b[9]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[9]) );
  DFFARX1 \add_combined_b_o_reg[8]  ( .D(add_combined_b[8]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[8]) );
  DFFARX1 \add_combined_b_o_reg[7]  ( .D(add_combined_b[7]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[7]) );
  DFFARX1 \add_combined_b_o_reg[6]  ( .D(add_combined_b[6]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[6]) );
  DFFARX1 \add_combined_b_o_reg[5]  ( .D(add_combined_b[5]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[5]) );
  DFFARX1 \add_combined_b_o_reg[4]  ( .D(add_combined_b[4]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[4]) );
  DFFARX1 \add_combined_b_o_reg[3]  ( .D(add_combined_b[3]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[3]) );
  DFFARX1 \add_combined_b_o_reg[2]  ( .D(add_combined_b[2]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[2]) );
  DFFARX1 \add_combined_b_o_reg[1]  ( .D(add_combined_b[1]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[1]) );
  DFFARX1 \add_combined_b_o_reg[0]  ( .D(add_combined_b[0]), .CLK(clk), .RSTB(
        n23), .Q(add_combined_b_o[0]) );
  DFFARX1 add_sign_a3_reg ( .D(add_sign_a2), .CLK(clk), .RSTB(n23), .Q(
        add_sign_a3) );
  AO22X1 U15 ( .IN1(N19), .IN2(n14), .IN3(n12), .IN4(N19), .Q(product[9]) );
  AO22X1 U16 ( .IN1(N18), .IN2(n20), .IN3(N18), .IN4(n11), .Q(product[8]) );
  AO22X1 U17 ( .IN1(N17), .IN2(n14), .IN3(N17), .IN4(n11), .Q(product[7]) );
  AO22X1 U18 ( .IN1(N16), .IN2(n14), .IN3(N16), .IN4(n11), .Q(product[6]) );
  AO22X1 U19 ( .IN1(N15), .IN2(n14), .IN3(N15), .IN4(n11), .Q(product[5]) );
  AND2X1 U20 ( .IN1(N60), .IN2(n11), .Q(product[50]) );
  AO22X1 U21 ( .IN1(N14), .IN2(n14), .IN3(N14), .IN4(n11), .Q(product[4]) );
  AND2X1 U22 ( .IN1(N59), .IN2(n13), .Q(product[49]) );
  AND2X1 U23 ( .IN1(N58), .IN2(n11), .Q(product[48]) );
  AND2X1 U24 ( .IN1(N57), .IN2(n12), .Q(product[47]) );
  AND2X1 U25 ( .IN1(N56), .IN2(n13), .Q(product[46]) );
  AND2X1 U26 ( .IN1(N55), .IN2(n13), .Q(product[45]) );
  AND2X1 U27 ( .IN1(N54), .IN2(n11), .Q(product[44]) );
  AND2X1 U28 ( .IN1(N53), .IN2(n12), .Q(product[43]) );
  AND2X1 U29 ( .IN1(N52), .IN2(n13), .Q(product[42]) );
  AND2X1 U30 ( .IN1(N51), .IN2(n11), .Q(product[41]) );
  AND2X1 U31 ( .IN1(N50), .IN2(n12), .Q(product[40]) );
  AO22X1 U32 ( .IN1(N13), .IN2(n14), .IN3(N13), .IN4(n12), .Q(product[3]) );
  AND2X1 U33 ( .IN1(N49), .IN2(n13), .Q(product[39]) );
  AND2X1 U34 ( .IN1(N48), .IN2(n13), .Q(product[38]) );
  AND2X1 U35 ( .IN1(N47), .IN2(n13), .Q(product[37]) );
  AND2X1 U36 ( .IN1(N46), .IN2(n13), .Q(product[36]) );
  AND2X1 U37 ( .IN1(N45), .IN2(n13), .Q(product[35]) );
  AND2X1 U38 ( .IN1(N44), .IN2(n13), .Q(product[34]) );
  AND2X1 U39 ( .IN1(N43), .IN2(n13), .Q(product[33]) );
  AND2X1 U40 ( .IN1(N42), .IN2(n13), .Q(product[32]) );
  AND2X1 U41 ( .IN1(N41), .IN2(n13), .Q(product[31]) );
  AND2X1 U42 ( .IN1(N40), .IN2(n13), .Q(product[30]) );
  AO22X1 U43 ( .IN1(N12), .IN2(n14), .IN3(N12), .IN4(n12), .Q(product[2]) );
  AND2X1 U44 ( .IN1(N39), .IN2(n13), .Q(product[29]) );
  AND2X1 U45 ( .IN1(N38), .IN2(n13), .Q(product[28]) );
  AND2X1 U46 ( .IN1(N37), .IN2(n12), .Q(product[27]) );
  AND2X1 U47 ( .IN1(N36), .IN2(n12), .Q(product[26]) );
  AO22X1 U49 ( .IN1(N34), .IN2(n14), .IN3(N34), .IN4(n12), .Q(product[24]) );
  AO22X1 U50 ( .IN1(N33), .IN2(n20), .IN3(N33), .IN4(n12), .Q(product[23]) );
  AO22X1 U51 ( .IN1(N32), .IN2(n20), .IN3(N32), .IN4(n12), .Q(product[22]) );
  AO22X1 U52 ( .IN1(N31), .IN2(n20), .IN3(N31), .IN4(n12), .Q(product[21]) );
  AO22X1 U53 ( .IN1(N30), .IN2(n20), .IN3(N30), .IN4(n12), .Q(product[20]) );
  AO22X1 U55 ( .IN1(N29), .IN2(n20), .IN3(N29), .IN4(n12), .Q(product[19]) );
  AO22X1 U56 ( .IN1(N28), .IN2(n20), .IN3(N28), .IN4(n12), .Q(product[18]) );
  AO22X1 U57 ( .IN1(N27), .IN2(n20), .IN3(N27), .IN4(n11), .Q(product[17]) );
  AO22X1 U58 ( .IN1(N26), .IN2(n14), .IN3(N26), .IN4(n11), .Q(product[16]) );
  AO22X1 U59 ( .IN1(N25), .IN2(n20), .IN3(N25), .IN4(n11), .Q(product[15]) );
  AO22X1 U60 ( .IN1(N24), .IN2(n14), .IN3(N24), .IN4(n11), .Q(product[14]) );
  AO22X1 U61 ( .IN1(N23), .IN2(n20), .IN3(N23), .IN4(n11), .Q(product[13]) );
  AO22X1 U62 ( .IN1(N22), .IN2(n14), .IN3(N22), .IN4(n11), .Q(product[12]) );
  AO22X1 U63 ( .IN1(N21), .IN2(n14), .IN3(N21), .IN4(n11), .Q(product[11]) );
  AO22X1 U64 ( .IN1(N20), .IN2(n14), .IN3(N20), .IN4(n12), .Q(product[10]) );
  AO22X1 U66 ( .IN1(add_exponent_a[7]), .IN2(n10), .IN3(N122), .IN4(n37), .Q(
        new_add_exponent[7]) );
  AO22X1 U67 ( .IN1(add_exponent_a[6]), .IN2(n15), .IN3(N121), .IN4(n8), .Q(
        new_add_exponent[6]) );
  AO22X1 U68 ( .IN1(add_exponent_a[5]), .IN2(n10), .IN3(N120), .IN4(n8), .Q(
        new_add_exponent[5]) );
  AO22X1 U69 ( .IN1(add_exponent_a[4]), .IN2(n10), .IN3(N119), .IN4(n8), .Q(
        new_add_exponent[4]) );
  AO22X1 U70 ( .IN1(add_exponent_a[3]), .IN2(n10), .IN3(N118), .IN4(n8), .Q(
        new_add_exponent[3]) );
  AO22X1 U71 ( .IN1(add_exponent_a[2]), .IN2(n15), .IN3(N117), .IN4(n8), .Q(
        new_add_exponent[2]) );
  AO22X1 U72 ( .IN1(add_exponent_a[1]), .IN2(n15), .IN3(N116), .IN4(n8), .Q(
        new_add_exponent[1]) );
  AO22X1 U73 ( .IN1(add_exponent_a[0]), .IN2(n15), .IN3(N115), .IN4(n8), .Q(
        new_add_exponent[0]) );
  AO22X1 U74 ( .IN1(N76), .IN2(n7), .IN3(add_fraction_b[9]), .IN4(n9), .Q(
        add_combined_b[9]) );
  AO22X1 U75 ( .IN1(N75), .IN2(n7), .IN3(add_fraction_b[8]), .IN4(n16), .Q(
        add_combined_b[8]) );
  AO22X1 U76 ( .IN1(N74), .IN2(n7), .IN3(add_fraction_b[7]), .IN4(n16), .Q(
        add_combined_b[7]) );
  AO22X1 U77 ( .IN1(N73), .IN2(n7), .IN3(add_fraction_b[6]), .IN4(n16), .Q(
        add_combined_b[6]) );
  AO22X1 U78 ( .IN1(N72), .IN2(n7), .IN3(add_fraction_b[5]), .IN4(n16), .Q(
        add_combined_b[5]) );
  AO22X1 U79 ( .IN1(N71), .IN2(n7), .IN3(add_fraction_b[4]), .IN4(n16), .Q(
        add_combined_b[4]) );
  AO22X1 U80 ( .IN1(N70), .IN2(n7), .IN3(add_fraction_b[3]), .IN4(n9), .Q(
        add_combined_b[3]) );
  AO22X1 U81 ( .IN1(N69), .IN2(n7), .IN3(add_fraction_b[2]), .IN4(n9), .Q(
        add_combined_b[2]) );
  AO21X1 U82 ( .IN1(N90), .IN2(n7), .IN3(n9), .Q(add_combined_b[23]) );
  AO22X1 U83 ( .IN1(N89), .IN2(n7), .IN3(add_fraction_b[22]), .IN4(n16), .Q(
        add_combined_b[22]) );
  AO22X1 U84 ( .IN1(N88), .IN2(n7), .IN3(add_fraction_b[21]), .IN4(n16), .Q(
        add_combined_b[21]) );
  AO22X1 U85 ( .IN1(N87), .IN2(n7), .IN3(add_fraction_b[20]), .IN4(n16), .Q(
        add_combined_b[20]) );
  AO22X1 U86 ( .IN1(N68), .IN2(n36), .IN3(add_fraction_b[1]), .IN4(n16), .Q(
        add_combined_b[1]) );
  AO22X1 U87 ( .IN1(N86), .IN2(n36), .IN3(add_fraction_b[19]), .IN4(n9), .Q(
        add_combined_b[19]) );
  AO22X1 U88 ( .IN1(N85), .IN2(n36), .IN3(add_fraction_b[18]), .IN4(n9), .Q(
        add_combined_b[18]) );
  AO22X1 U89 ( .IN1(N84), .IN2(n7), .IN3(add_fraction_b[17]), .IN4(n9), .Q(
        add_combined_b[17]) );
  AO22X1 U90 ( .IN1(N83), .IN2(n7), .IN3(add_fraction_b[16]), .IN4(n9), .Q(
        add_combined_b[16]) );
  AO22X1 U91 ( .IN1(N82), .IN2(n36), .IN3(add_fraction_b[15]), .IN4(n9), .Q(
        add_combined_b[15]) );
  AO22X1 U92 ( .IN1(N81), .IN2(n36), .IN3(add_fraction_b[14]), .IN4(n9), .Q(
        add_combined_b[14]) );
  AO22X1 U93 ( .IN1(N80), .IN2(n36), .IN3(add_fraction_b[13]), .IN4(n9), .Q(
        add_combined_b[13]) );
  AO22X1 U94 ( .IN1(N79), .IN2(n36), .IN3(add_fraction_b[12]), .IN4(n9), .Q(
        add_combined_b[12]) );
  AO22X1 U95 ( .IN1(N78), .IN2(n36), .IN3(add_fraction_b[11]), .IN4(n9), .Q(
        add_combined_b[11]) );
  AO22X1 U96 ( .IN1(N77), .IN2(n36), .IN3(add_fraction_b[10]), .IN4(n9), .Q(
        add_combined_b[10]) );
  AO22X1 U97 ( .IN1(N67), .IN2(n7), .IN3(add_fraction_b[0]), .IN4(n9), .Q(
        add_combined_b[0]) );
  AO22X1 U98 ( .IN1(add_fraction_a[9]), .IN2(n15), .IN3(N100), .IN4(n8), .Q(
        add_combined_a[9]) );
  AO22X1 U99 ( .IN1(add_fraction_a[8]), .IN2(n15), .IN3(N99), .IN4(n8), .Q(
        add_combined_a[8]) );
  AO22X1 U100 ( .IN1(add_fraction_a[7]), .IN2(n15), .IN3(N98), .IN4(n8), .Q(
        add_combined_a[7]) );
  AO22X1 U101 ( .IN1(add_fraction_a[6]), .IN2(n15), .IN3(N97), .IN4(n8), .Q(
        add_combined_a[6]) );
  AO22X1 U102 ( .IN1(add_fraction_a[5]), .IN2(n15), .IN3(N96), .IN4(n37), .Q(
        add_combined_a[5]) );
  AO22X1 U103 ( .IN1(add_fraction_a[4]), .IN2(n15), .IN3(N95), .IN4(n37), .Q(
        add_combined_a[4]) );
  AO22X1 U104 ( .IN1(add_fraction_a[3]), .IN2(n15), .IN3(N94), .IN4(n37), .Q(
        add_combined_a[3]) );
  AO22X1 U105 ( .IN1(add_fraction_a[2]), .IN2(n15), .IN3(N93), .IN4(n37), .Q(
        add_combined_a[2]) );
  AO21X1 U106 ( .IN1(N114), .IN2(n8), .IN3(n10), .Q(add_combined_a[23]) );
  AO22X1 U107 ( .IN1(add_fraction_a[22]), .IN2(n10), .IN3(N113), .IN4(n37), 
        .Q(add_combined_a[22]) );
  AO22X1 U108 ( .IN1(add_fraction_a[21]), .IN2(n10), .IN3(N112), .IN4(n37), 
        .Q(add_combined_a[21]) );
  AO22X1 U109 ( .IN1(add_fraction_a[20]), .IN2(n10), .IN3(N111), .IN4(n37), 
        .Q(add_combined_a[20]) );
  AO22X1 U110 ( .IN1(add_fraction_a[1]), .IN2(n10), .IN3(N92), .IN4(n37), .Q(
        add_combined_a[1]) );
  AO22X1 U111 ( .IN1(add_fraction_a[19]), .IN2(n10), .IN3(N110), .IN4(n37), 
        .Q(add_combined_a[19]) );
  AO22X1 U112 ( .IN1(add_fraction_a[18]), .IN2(n15), .IN3(N109), .IN4(n37), 
        .Q(add_combined_a[18]) );
  AO22X1 U113 ( .IN1(add_fraction_a[17]), .IN2(n10), .IN3(N108), .IN4(n37), 
        .Q(add_combined_a[17]) );
  AO22X1 U114 ( .IN1(add_fraction_a[16]), .IN2(n10), .IN3(N107), .IN4(n37), 
        .Q(add_combined_a[16]) );
  AO22X1 U115 ( .IN1(add_fraction_a[15]), .IN2(n10), .IN3(N106), .IN4(n37), 
        .Q(add_combined_a[15]) );
  AO22X1 U116 ( .IN1(add_fraction_a[14]), .IN2(n10), .IN3(N105), .IN4(n37), 
        .Q(add_combined_a[14]) );
  AO22X1 U117 ( .IN1(add_fraction_a[13]), .IN2(n10), .IN3(N104), .IN4(n37), 
        .Q(add_combined_a[13]) );
  AO22X1 U118 ( .IN1(add_fraction_a[12]), .IN2(n10), .IN3(N103), .IN4(n37), 
        .Q(add_combined_a[12]) );
  AO22X1 U119 ( .IN1(add_fraction_a[11]), .IN2(n10), .IN3(N102), .IN4(n8), .Q(
        add_combined_a[11]) );
  AO22X1 U120 ( .IN1(add_fraction_a[10]), .IN2(n10), .IN3(N101), .IN4(n37), 
        .Q(add_combined_a[10]) );
  AO22X1 U121 ( .IN1(add_fraction_a[0]), .IN2(n15), .IN3(N91), .IN4(n8), .Q(
        add_combined_a[0]) );
  NAND3X0 U122 ( .IN1(n39), .IN2(n38), .IN3(add_lesser_flag), .QN(n17) );
  NAND3X0 U123 ( .IN1(n39), .IN2(n40), .IN3(add_zero_flag), .QN(n18) );
  NAND3X0 U124 ( .IN1(n40), .IN2(n38), .IN3(add_greater_flag), .QN(n19) );
  booth_DW01_add_0 add_128 ( .A(add_exponent_a), .B({add_difference[7:3], n6, 
        add_difference[1:0]}), .CI(1'b0), .SUM({N122, N121, N120, N119, N118, 
        N117, N116, N115}) );
  booth_DW_rash_0 srl_127 ( .A({1'b1, add_fraction_a}), .DATA_TC(1'b0), .SH({
        add_difference[7:3], n6, n4, add_difference[0]}), .SH_TC(1'b0), .B({
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91}) );
  booth_DW_rash_1 srl_118 ( .A({1'b1, add_fraction_b}), .DATA_TC(1'b0), .SH({
        add_difference[7:3], n6, n4, add_difference[0]}), .SH_TC(1'b0), .B({
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, N74, N73, N72, N71, N70, N69, N68, N67}) );
  NAND2X1 U3 ( .IN1(n19), .IN2(n18), .QN(n10) );
  NBUFFX2 U4 ( .INP(add_difference[1]), .Z(n4) );
  NBUFFX2 U5 ( .INP(n16), .Z(n9) );
  NBUFFX2 U6 ( .INP(n37), .Z(n8) );
  NBUFFX2 U7 ( .INP(n36), .Z(n7) );
  NBUFFX2 U8 ( .INP(n21), .Z(n23) );
  NBUFFX2 U12 ( .INP(n21), .Z(n24) );
  NBUFFX2 U13 ( .INP(n21), .Z(n25) );
  NBUFFX2 U14 ( .INP(n21), .Z(n26) );
  NBUFFX2 U48 ( .INP(n21), .Z(n27) );
  NBUFFX2 U54 ( .INP(n21), .Z(n28) );
  NBUFFX2 U65 ( .INP(n21), .Z(n29) );
  NBUFFX2 U125 ( .INP(n21), .Z(n31) );
  NBUFFX2 U126 ( .INP(n22), .Z(n33) );
  NBUFFX2 U127 ( .INP(n22), .Z(n34) );
  NBUFFX2 U128 ( .INP(n21), .Z(n30) );
  NBUFFX2 U129 ( .INP(n21), .Z(n32) );
  NBUFFX2 U130 ( .INP(n22), .Z(n35) );
  NAND2X1 U131 ( .IN1(n19), .IN2(n18), .QN(n15) );
  INVX0 U132 ( .INP(n17), .ZN(n37) );
  NAND2X1 U133 ( .IN1(n17), .IN2(n18), .QN(n16) );
  INVX0 U134 ( .INP(n19), .ZN(n36) );
  NBUFFX2 U135 ( .INP(reset), .Z(n21) );
  NBUFFX2 U136 ( .INP(reset), .Z(n22) );
  INVX0 U137 ( .INP(combined_a[0]), .ZN(n20) );
  INVX0 U138 ( .INP(combined_a[0]), .ZN(n14) );
  INVX0 U139 ( .INP(add_greater_flag), .ZN(n39) );
  INVX0 U140 ( .INP(add_zero_flag), .ZN(n38) );
  INVX0 U141 ( .INP(add_lesser_flag), .ZN(n40) );
  INVX0 U143 ( .INP(add_difference[2]), .ZN(n5) );
  INVX0 U144 ( .INP(n5), .ZN(n6) );
  INVX0 U145 ( .INP(n20), .ZN(n11) );
  INVX0 U146 ( .INP(n20), .ZN(n12) );
  INVX0 U147 ( .INP(n14), .ZN(n13) );
endmodule


module booth2_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51;
  wire   [25:0] carry;

  FADDX1 U2_23 ( .A(A[23]), .B(n28), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n29), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n34), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n39), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_1 ( .A(A[1]), .B(n50), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  FADDX1 U2_11 ( .A(A[11]), .B(n40), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n42), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n45), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_21 ( .A(A[21]), .B(n30), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n33), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n36), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n46), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n49), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_16 ( .A(A[16]), .B(n35), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n38), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n37), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  NAND2X0 U1 ( .IN1(A[19]), .IN2(carry[19]), .QN(n2) );
  XOR3X1 U2 ( .IN1(A[19]), .IN2(n32), .IN3(carry[19]), .Q(DIFF[19]) );
  NAND2X1 U3 ( .IN1(A[19]), .IN2(n32), .QN(n1) );
  NAND2X0 U4 ( .IN1(n32), .IN2(carry[19]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[20]) );
  XOR2X1 U6 ( .IN1(A[20]), .IN2(n31), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[20]), .Q(DIFF[20]) );
  NAND2X0 U8 ( .IN1(A[20]), .IN2(n31), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[20]), .IN2(carry[20]), .QN(n6) );
  NAND2X0 U10 ( .IN1(n31), .IN2(carry[20]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[21]) );
  INVX0 U12 ( .INP(B[10]), .ZN(n41) );
  XNOR2X1 U13 ( .IN1(n8), .IN2(carry[8]), .Q(DIFF[8]) );
  XNOR2X1 U14 ( .IN1(A[8]), .IN2(n43), .Q(n8) );
  XOR3X2 U15 ( .IN1(A[7]), .IN2(n44), .IN3(carry[7]), .Q(DIFF[7]) );
  NAND2X0 U16 ( .IN1(A[7]), .IN2(n44), .QN(n9) );
  NAND2X0 U17 ( .IN1(A[7]), .IN2(carry[7]), .QN(n10) );
  NAND2X0 U18 ( .IN1(n44), .IN2(carry[7]), .QN(n11) );
  NAND3X0 U19 ( .IN1(n9), .IN2(n10), .IN3(n11), .QN(carry[8]) );
  NAND2X0 U20 ( .IN1(A[8]), .IN2(n43), .QN(n12) );
  NAND2X0 U21 ( .IN1(A[8]), .IN2(carry[8]), .QN(n13) );
  NAND2X0 U22 ( .IN1(n43), .IN2(carry[8]), .QN(n14) );
  NAND3X0 U23 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[9]) );
  XOR3X1 U24 ( .IN1(A[3]), .IN2(n48), .IN3(carry[3]), .Q(DIFF[3]) );
  NAND2X1 U25 ( .IN1(A[3]), .IN2(n48), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[3]), .IN2(carry[3]), .QN(n16) );
  NAND2X0 U27 ( .IN1(n48), .IN2(carry[3]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[4]) );
  XOR2X1 U29 ( .IN1(A[4]), .IN2(n47), .Q(n18) );
  XOR2X1 U30 ( .IN1(n18), .IN2(carry[4]), .Q(DIFF[4]) );
  NAND2X0 U31 ( .IN1(A[4]), .IN2(n47), .QN(n19) );
  NAND2X0 U32 ( .IN1(A[4]), .IN2(carry[4]), .QN(n20) );
  NAND2X0 U33 ( .IN1(n47), .IN2(carry[4]), .QN(n21) );
  NAND3X0 U34 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[5]) );
  XOR3X1 U35 ( .IN1(carry[10]), .IN2(n41), .IN3(A[10]), .Q(DIFF[10]) );
  NAND2X0 U36 ( .IN1(A[10]), .IN2(carry[10]), .QN(n22) );
  NAND2X0 U37 ( .IN1(n41), .IN2(carry[10]), .QN(n23) );
  NAND2X0 U38 ( .IN1(n41), .IN2(A[10]), .QN(n24) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n24), .IN3(n23), .QN(carry[11]) );
  NAND2X0 U40 ( .IN1(n25), .IN2(n26), .QN(carry[1]) );
  INVX0 U41 ( .INP(carry[24]), .ZN(DIFF[24]) );
  INVX0 U42 ( .INP(B[1]), .ZN(n50) );
  INVX0 U43 ( .INP(A[0]), .ZN(n25) );
  INVX0 U44 ( .INP(n51), .ZN(n26) );
  INVX0 U45 ( .INP(B[0]), .ZN(n51) );
  INVX0 U46 ( .INP(B[13]), .ZN(n38) );
  INVX0 U47 ( .INP(B[14]), .ZN(n37) );
  INVX0 U48 ( .INP(B[15]), .ZN(n36) );
  INVX0 U49 ( .INP(B[16]), .ZN(n35) );
  INVX0 U50 ( .INP(B[17]), .ZN(n34) );
  INVX0 U51 ( .INP(B[18]), .ZN(n33) );
  INVX0 U52 ( .INP(B[19]), .ZN(n32) );
  INVX0 U53 ( .INP(B[12]), .ZN(n39) );
  INVX0 U54 ( .INP(B[20]), .ZN(n31) );
  INVX0 U55 ( .INP(B[11]), .ZN(n40) );
  INVX0 U56 ( .INP(B[21]), .ZN(n30) );
  INVX0 U57 ( .INP(B[22]), .ZN(n29) );
  INVX0 U58 ( .INP(B[9]), .ZN(n42) );
  INVX0 U59 ( .INP(B[3]), .ZN(n48) );
  INVX0 U60 ( .INP(B[4]), .ZN(n47) );
  INVX0 U61 ( .INP(B[5]), .ZN(n46) );
  INVX0 U62 ( .INP(B[6]), .ZN(n45) );
  INVX0 U63 ( .INP(B[7]), .ZN(n44) );
  INVX0 U64 ( .INP(B[8]), .ZN(n43) );
  INVX0 U65 ( .INP(B[23]), .ZN(n28) );
  XOR2X1 U66 ( .IN1(n26), .IN2(A[0]), .Q(DIFF[0]) );
  INVX0 U67 ( .INP(B[2]), .ZN(n49) );
endmodule


module booth2_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47;
  wire   [25:0] carry;

  FADDX1 U2_16 ( .A(A[16]), .B(n31), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n25), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n28), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n42), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_17 ( .A(A[17]), .B(n30), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n33), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_11 ( .A(n20), .B(n36), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n41), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n44), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_18 ( .A(A[18]), .B(n29), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n32), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n35), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_8 ( .A(A[8]), .B(n39), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n43), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n46), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  FADDX1 U2_13 ( .A(A[13]), .B(n34), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n40), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n45), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  INVX0 U1 ( .INP(B[23]), .ZN(n24) );
  XOR3X1 U2 ( .IN1(A[20]), .IN2(n27), .IN3(carry[20]), .Q(DIFF[20]) );
  XOR2X1 U3 ( .IN1(n24), .IN2(A[23]), .Q(n8) );
  AND3X1 U4 ( .IN1(n9), .IN2(n11), .IN3(n10), .Q(DIFF[24]) );
  XOR3X1 U5 ( .IN1(A[9]), .IN2(n38), .IN3(carry[9]), .Q(DIFF[9]) );
  NAND2X1 U6 ( .IN1(A[9]), .IN2(n38), .QN(n1) );
  NAND2X1 U7 ( .IN1(A[9]), .IN2(carry[9]), .QN(n2) );
  NAND2X0 U8 ( .IN1(n38), .IN2(carry[9]), .QN(n3) );
  NAND3X0 U9 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[10]) );
  XOR2X1 U10 ( .IN1(A[10]), .IN2(n37), .Q(n4) );
  XOR2X1 U11 ( .IN1(n4), .IN2(carry[10]), .Q(DIFF[10]) );
  NAND2X0 U12 ( .IN1(A[10]), .IN2(n37), .QN(n5) );
  NAND2X0 U13 ( .IN1(A[10]), .IN2(carry[10]), .QN(n6) );
  NAND2X0 U14 ( .IN1(n37), .IN2(carry[10]), .QN(n7) );
  NAND3X0 U15 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[11]) );
  XOR2X1 U16 ( .IN1(n8), .IN2(carry[23]), .Q(DIFF[23]) );
  NAND2X0 U17 ( .IN1(A[23]), .IN2(carry[23]), .QN(n9) );
  NAND2X0 U18 ( .IN1(n24), .IN2(carry[23]), .QN(n10) );
  NAND2X0 U19 ( .IN1(n24), .IN2(A[23]), .QN(n11) );
  NAND2X0 U20 ( .IN1(A[20]), .IN2(n27), .QN(n12) );
  NAND2X0 U21 ( .IN1(A[20]), .IN2(carry[20]), .QN(n13) );
  NAND2X0 U22 ( .IN1(n27), .IN2(carry[20]), .QN(n14) );
  NAND3X0 U23 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[21]) );
  XOR2X1 U24 ( .IN1(A[21]), .IN2(n26), .Q(n15) );
  XOR2X1 U25 ( .IN1(n15), .IN2(carry[21]), .Q(DIFF[21]) );
  NAND2X0 U26 ( .IN1(A[21]), .IN2(n26), .QN(n16) );
  NAND2X0 U27 ( .IN1(A[21]), .IN2(carry[21]), .QN(n17) );
  NAND2X0 U28 ( .IN1(n26), .IN2(carry[21]), .QN(n18) );
  NAND3X0 U29 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[22]) );
  INVX0 U30 ( .INP(A[11]), .ZN(n19) );
  INVX0 U31 ( .INP(n19), .ZN(n20) );
  NAND2X0 U32 ( .IN1(n21), .IN2(n22), .QN(carry[1]) );
  INVX0 U33 ( .INP(A[0]), .ZN(n21) );
  INVX0 U34 ( .INP(B[14]), .ZN(n33) );
  INVX0 U35 ( .INP(B[16]), .ZN(n31) );
  INVX0 U36 ( .INP(B[8]), .ZN(n39) );
  INVX0 U37 ( .INP(B[4]), .ZN(n43) );
  INVX0 U38 ( .INP(B[6]), .ZN(n41) );
  INVX0 U39 ( .INP(B[18]), .ZN(n29) );
  INVX0 U40 ( .INP(B[12]), .ZN(n35) );
  INVX0 U41 ( .INP(B[20]), .ZN(n27) );
  INVX0 U42 ( .INP(B[9]), .ZN(n38) );
  INVX0 U43 ( .INP(B[10]), .ZN(n37) );
  INVX0 U44 ( .INP(B[13]), .ZN(n34) );
  INVX0 U45 ( .INP(B[15]), .ZN(n32) );
  INVX0 U46 ( .INP(B[17]), .ZN(n30) );
  INVX0 U47 ( .INP(B[19]), .ZN(n28) );
  INVX0 U48 ( .INP(B[11]), .ZN(n36) );
  INVX0 U49 ( .INP(B[21]), .ZN(n26) );
  INVX0 U50 ( .INP(B[22]), .ZN(n25) );
  INVX0 U51 ( .INP(B[3]), .ZN(n44) );
  INVX0 U52 ( .INP(B[7]), .ZN(n40) );
  INVX0 U53 ( .INP(B[5]), .ZN(n42) );
  INVX0 U54 ( .INP(n47), .ZN(n22) );
  XOR2X1 U55 ( .IN1(n22), .IN2(A[0]), .Q(DIFF[0]) );
  INVX0 U56 ( .INP(B[2]), .ZN(n45) );
  INVX0 U57 ( .INP(B[1]), .ZN(n46) );
  INVX0 U58 ( .INP(B[0]), .ZN(n47) );
endmodule


module booth2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n23), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X1 U2 ( .IN1(A[46]), .IN2(B[46]), .QN(n1) );
  NAND2X1 U3 ( .IN1(A[46]), .IN2(carry[46]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[46]), .IN2(carry[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[47]) );
  XOR2X1 U6 ( .IN1(A[47]), .IN2(B[47]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[47]), .Q(SUM[47]) );
  NAND2X0 U8 ( .IN1(A[47]), .IN2(B[47]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[47]), .IN2(carry[47]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[47]), .IN2(carry[47]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[48]) );
  XOR3X2 U12 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U13 ( .IN1(A[38]), .IN2(B[38]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[38]), .IN2(carry[38]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[38]), .IN2(carry[38]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[39]) );
  XOR2X1 U17 ( .IN1(A[39]), .IN2(B[39]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U19 ( .IN1(A[39]), .IN2(B[39]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[39]), .IN2(carry[39]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[39]), .IN2(carry[39]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[40]) );
  DELLN2X2 U23 ( .INP(carry[41]), .Z(n15) );
  XOR3X2 U24 ( .IN1(carry[40]), .IN2(B[40]), .IN3(A[40]), .Q(SUM[40]) );
  NAND2X0 U25 ( .IN1(A[40]), .IN2(B[40]), .QN(n16) );
  NAND2X0 U26 ( .IN1(A[40]), .IN2(carry[40]), .QN(n17) );
  NAND2X0 U27 ( .IN1(B[40]), .IN2(carry[40]), .QN(n18) );
  NAND3X0 U28 ( .IN1(n17), .IN2(n18), .IN3(n16), .QN(carry[41]) );
  XOR2X1 U29 ( .IN1(A[41]), .IN2(B[41]), .Q(n19) );
  XOR2X1 U30 ( .IN1(n19), .IN2(n15), .Q(SUM[41]) );
  NAND2X0 U31 ( .IN1(A[41]), .IN2(B[41]), .QN(n20) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(carry[41]), .QN(n21) );
  NAND2X0 U33 ( .IN1(B[41]), .IN2(carry[41]), .QN(n22) );
  NAND3X0 U34 ( .IN1(n21), .IN2(n22), .IN3(n20), .QN(carry[42]) );
  AND2X1 U35 ( .IN1(A[26]), .IN2(B[26]), .Q(n23) );
  XOR2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n26), .CO(carry[28]), .S(SUM[27])
         );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX2 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX2 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  XOR2X1 U1 ( .IN1(A[50]), .IN2(carry[50]), .Q(SUM[50]) );
  XOR3X1 U2 ( .IN1(carry[43]), .IN2(B[43]), .IN3(A[43]), .Q(SUM[43]) );
  NAND2X1 U3 ( .IN1(A[43]), .IN2(carry[43]), .QN(n1) );
  NAND2X0 U4 ( .IN1(B[43]), .IN2(carry[43]), .QN(n2) );
  NAND2X1 U5 ( .IN1(B[43]), .IN2(A[43]), .QN(n3) );
  NAND3X0 U6 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[44]) );
  XOR3X1 U7 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U8 ( .IN1(A[41]), .IN2(B[41]), .IN3(carry[41]), .Q(SUM[41]) );
  NAND2X1 U9 ( .IN1(A[41]), .IN2(B[41]), .QN(n4) );
  NAND2X1 U10 ( .IN1(A[41]), .IN2(carry[41]), .QN(n5) );
  NAND2X0 U11 ( .IN1(B[41]), .IN2(carry[41]), .QN(n6) );
  NAND3X0 U12 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[42]) );
  XOR2X1 U13 ( .IN1(A[42]), .IN2(B[42]), .Q(n7) );
  XOR2X1 U14 ( .IN1(n7), .IN2(carry[42]), .Q(SUM[42]) );
  NAND2X0 U15 ( .IN1(A[42]), .IN2(B[42]), .QN(n8) );
  NAND2X0 U16 ( .IN1(A[42]), .IN2(carry[42]), .QN(n9) );
  NAND2X0 U17 ( .IN1(B[42]), .IN2(carry[42]), .QN(n10) );
  NAND3X0 U18 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[43]) );
  XOR2X1 U19 ( .IN1(n22), .IN2(carry[48]), .Q(SUM[48]) );
  DELLN2X2 U20 ( .INP(carry[45]), .Z(n11) );
  XOR3X2 U21 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U22 ( .IN1(A[44]), .IN2(B[44]), .QN(n12) );
  NAND2X0 U23 ( .IN1(A[44]), .IN2(carry[44]), .QN(n13) );
  NAND2X0 U24 ( .IN1(B[44]), .IN2(carry[44]), .QN(n14) );
  NAND3X0 U25 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[45]) );
  XOR2X1 U26 ( .IN1(A[45]), .IN2(B[45]), .Q(n15) );
  XOR2X1 U27 ( .IN1(n15), .IN2(n11), .Q(SUM[45]) );
  NAND2X0 U28 ( .IN1(A[45]), .IN2(B[45]), .QN(n16) );
  NAND2X0 U29 ( .IN1(A[45]), .IN2(carry[45]), .QN(n17) );
  NAND2X0 U30 ( .IN1(B[45]), .IN2(carry[45]), .QN(n18) );
  NAND3X0 U31 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[46]) );
  NAND2X0 U32 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U33 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U34 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U35 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[48]) );
  XOR2X1 U36 ( .IN1(A[48]), .IN2(B[48]), .Q(n22) );
  NAND2X0 U37 ( .IN1(A[48]), .IN2(B[48]), .QN(n23) );
  NAND2X0 U38 ( .IN1(A[48]), .IN2(carry[48]), .QN(n24) );
  NAND2X0 U39 ( .IN1(B[48]), .IN2(carry[48]), .QN(n25) );
  NAND3X0 U40 ( .IN1(n23), .IN2(n24), .IN3(n25), .QN(carry[49]) );
  AND2X1 U41 ( .IN1(A[26]), .IN2(B[26]), .Q(n26) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth2_DW01_add_2 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [24:1] carry;

  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n26), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_11 ( .A(n7), .B(carry[11]), .CI(B[11]), .CO(carry[12]), .S(SUM[11]) );
  INVX0 U1 ( .INP(carry[22]), .ZN(n1) );
  INVX0 U2 ( .INP(n1), .ZN(n2) );
  XOR3X1 U3 ( .IN1(carry[10]), .IN2(B[10]), .IN3(A[10]), .Q(SUM[10]) );
  NAND2X1 U4 ( .IN1(A[10]), .IN2(carry[10]), .QN(n3) );
  NAND2X0 U5 ( .IN1(B[10]), .IN2(carry[10]), .QN(n4) );
  NAND2X0 U6 ( .IN1(B[10]), .IN2(A[10]), .QN(n5) );
  NAND3X0 U7 ( .IN1(n3), .IN2(n5), .IN3(n4), .QN(carry[11]) );
  INVX0 U8 ( .INP(A[11]), .ZN(n6) );
  INVX0 U9 ( .INP(n6), .ZN(n7) );
  XOR3X1 U10 ( .IN1(n2), .IN2(A[22]), .IN3(B[22]), .Q(SUM[22]) );
  NAND2X0 U11 ( .IN1(B[22]), .IN2(carry[22]), .QN(n8) );
  NAND2X0 U12 ( .IN1(A[22]), .IN2(carry[22]), .QN(n9) );
  NAND2X0 U13 ( .IN1(A[22]), .IN2(B[22]), .QN(n10) );
  NAND3X0 U14 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[23]) );
  DELLN2X2 U15 ( .INP(carry[21]), .Z(n11) );
  XOR3X1 U16 ( .IN1(A[20]), .IN2(B[20]), .IN3(carry[20]), .Q(SUM[20]) );
  XNOR2X1 U17 ( .IN1(n12), .IN2(carry[7]), .Q(SUM[7]) );
  XNOR2X1 U18 ( .IN1(A[7]), .IN2(B[7]), .Q(n12) );
  XOR3X1 U19 ( .IN1(A[6]), .IN2(B[6]), .IN3(carry[6]), .Q(SUM[6]) );
  NAND2X0 U20 ( .IN1(A[6]), .IN2(B[6]), .QN(n13) );
  NAND2X0 U21 ( .IN1(A[6]), .IN2(carry[6]), .QN(n14) );
  NAND2X0 U22 ( .IN1(B[6]), .IN2(carry[6]), .QN(n15) );
  NAND3X0 U23 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[7]) );
  NAND2X0 U24 ( .IN1(A[7]), .IN2(B[7]), .QN(n16) );
  NAND2X0 U25 ( .IN1(A[7]), .IN2(carry[7]), .QN(n17) );
  NAND2X0 U26 ( .IN1(B[7]), .IN2(carry[7]), .QN(n18) );
  NAND3X0 U27 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[8]) );
  NAND2X0 U28 ( .IN1(A[20]), .IN2(B[20]), .QN(n19) );
  NAND2X0 U29 ( .IN1(A[20]), .IN2(carry[20]), .QN(n20) );
  NAND2X0 U30 ( .IN1(B[20]), .IN2(carry[20]), .QN(n21) );
  NAND3X0 U31 ( .IN1(n21), .IN2(n20), .IN3(n19), .QN(carry[21]) );
  XOR2X1 U32 ( .IN1(A[21]), .IN2(B[21]), .Q(n22) );
  XOR2X1 U33 ( .IN1(n22), .IN2(n11), .Q(SUM[21]) );
  NAND2X0 U34 ( .IN1(A[21]), .IN2(B[21]), .QN(n23) );
  NAND2X0 U35 ( .IN1(A[21]), .IN2(carry[21]), .QN(n24) );
  NAND2X0 U36 ( .IN1(B[21]), .IN2(carry[21]), .QN(n25) );
  NAND3X0 U37 ( .IN1(n25), .IN2(n24), .IN3(n23), .QN(carry[22]) );
  AND2X1 U38 ( .IN1(A[0]), .IN2(B[0]), .Q(n26) );
  XOR2X1 U39 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module booth2 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_sign_a, add_sign_b, add_new_a, 
        add_new_b, add_sum_o, add_new_add_sign_o, add_sign_a3, add_sign_b3, 
        add_new_exponent, add_new_exponent2, s, s2, add_greater_flag2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [23:0] add_new_a;
  input [23:0] add_new_b;
  output [24:0] add_sum_o;
  input [7:0] add_new_exponent;
  output [7:0] add_new_exponent2;
  input clk, reset, new_sign, add_sign_a, add_sign_b, s, add_greater_flag2;
  output new_sign2, add_new_add_sign_o, add_sign_a3, add_sign_b3, s2;
  wire   N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, add_new_sign, N124, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, n16, n17, n18, n19, n22, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n20, n21, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   [24:0] add_sum;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[24] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n117), .Q(new_sign2)
         );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n117), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n117), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n116), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n115), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n114), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n113), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n112), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(1'b0), .CLK(clk), .RSTB(n112), .Q(
        combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n112), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n111), 
        .Q(combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n20), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n29), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n37), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n44), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n50), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n58), .CLK(clk), .RSTB(n111), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n68), .CLK(clk), .RSTB(n110), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n110), 
        .Q(combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n110), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n109), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n109), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n109), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n109), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n109), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n109), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n11), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n24), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n32), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n40), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n46), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n53), .CLK(clk), .RSTB(n109), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n62), .CLK(clk), .RSTB(n108), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n73), .CLK(clk), .RSTB(n108), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n108), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n108), 
        .Q(new_exponent2[0]) );
  DFFARX1 add_sign_b3_reg ( .D(add_sign_b), .CLK(clk), .RSTB(n107), .Q(
        add_sign_b3) );
  DFFARX1 \add_new_exponent2_reg[7]  ( .D(add_new_exponent[7]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[7]) );
  DFFARX1 \add_new_exponent2_reg[6]  ( .D(add_new_exponent[6]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[6]) );
  DFFARX1 \add_new_exponent2_reg[5]  ( .D(add_new_exponent[5]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[5]) );
  DFFARX1 \add_new_exponent2_reg[4]  ( .D(add_new_exponent[4]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[4]) );
  DFFARX1 \add_new_exponent2_reg[3]  ( .D(add_new_exponent[3]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[3]) );
  DFFARX1 \add_new_exponent2_reg[2]  ( .D(add_new_exponent[2]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[2]) );
  DFFARX1 \add_new_exponent2_reg[1]  ( .D(add_new_exponent[1]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[1]) );
  DFFARX1 \add_new_exponent2_reg[0]  ( .D(add_new_exponent[0]), .CLK(clk), 
        .RSTB(n107), .Q(add_new_exponent2[0]) );
  DFFARX1 add_new_add_sign_o_reg ( .D(add_new_sign), .CLK(clk), .RSTB(n107), 
        .Q(add_new_add_sign_o) );
  DFFARX1 \add_sum_o_reg[24]  ( .D(add_sum[24]), .CLK(clk), .RSTB(n107), .Q(
        add_sum_o[24]) );
  DFFARX1 \add_sum_o_reg[23]  ( .D(add_sum[23]), .CLK(clk), .RSTB(n107), .Q(
        add_sum_o[23]) );
  DFFARX1 \add_sum_o_reg[22]  ( .D(add_sum[22]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[22]) );
  DFFARX1 \add_sum_o_reg[21]  ( .D(add_sum[21]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[21]) );
  DFFARX1 \add_sum_o_reg[20]  ( .D(add_sum[20]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[20]) );
  DFFARX1 \add_sum_o_reg[19]  ( .D(add_sum[19]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[19]) );
  DFFARX1 \add_sum_o_reg[18]  ( .D(add_sum[18]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[18]) );
  DFFARX1 \add_sum_o_reg[17]  ( .D(add_sum[17]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[17]) );
  DFFARX1 \add_sum_o_reg[16]  ( .D(add_sum[16]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[16]) );
  DFFARX1 \add_sum_o_reg[15]  ( .D(add_sum[15]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[15]) );
  DFFARX1 \add_sum_o_reg[14]  ( .D(add_sum[14]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[14]) );
  DFFARX1 \add_sum_o_reg[13]  ( .D(add_sum[13]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[13]) );
  DFFARX1 \add_sum_o_reg[12]  ( .D(add_sum[12]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[12]) );
  DFFARX1 \add_sum_o_reg[11]  ( .D(add_sum[11]), .CLK(clk), .RSTB(n106), .Q(
        add_sum_o[11]) );
  DFFARX1 \add_sum_o_reg[10]  ( .D(add_sum[10]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[10]) );
  DFFARX1 \add_sum_o_reg[9]  ( .D(add_sum[9]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[9]) );
  DFFARX1 \add_sum_o_reg[8]  ( .D(add_sum[8]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[8]) );
  DFFARX1 \add_sum_o_reg[7]  ( .D(add_sum[7]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[7]) );
  DFFARX1 \add_sum_o_reg[6]  ( .D(add_sum[6]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[6]) );
  DFFARX1 \add_sum_o_reg[5]  ( .D(add_sum[5]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[5]) );
  DFFARX1 \add_sum_o_reg[4]  ( .D(add_sum[4]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[4]) );
  DFFARX1 \add_sum_o_reg[3]  ( .D(add_sum[3]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[3]) );
  DFFARX1 \add_sum_o_reg[2]  ( .D(add_sum[2]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[2]) );
  DFFARX1 \add_sum_o_reg[1]  ( .D(add_sum[1]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[1]) );
  DFFARX1 \add_sum_o_reg[0]  ( .D(add_sum[0]), .CLK(clk), .RSTB(n105), .Q(
        add_sum_o[0]) );
  DFFARX1 add_sign_a3_reg ( .D(add_sign_a), .CLK(clk), .RSTB(n105), .Q(
        add_sign_a3) );
  AO222X1 U13 ( .IN1(N29), .IN2(n100), .IN3(N80), .IN4(n97), .IN5(
        product_shift[9]), .IN6(n95), .Q(product2[9]) );
  AO222X1 U14 ( .IN1(N28), .IN2(n100), .IN3(N79), .IN4(n97), .IN5(
        product_shift[8]), .IN6(n18), .Q(product2[8]) );
  AO222X1 U15 ( .IN1(N27), .IN2(n100), .IN3(N78), .IN4(n97), .IN5(
        product_shift[7]), .IN6(n18), .Q(product2[7]) );
  AO222X1 U16 ( .IN1(N26), .IN2(n100), .IN3(N77), .IN4(n97), .IN5(
        product_shift[6]), .IN6(n18), .Q(product2[6]) );
  AO222X1 U17 ( .IN1(N25), .IN2(n100), .IN3(N76), .IN4(n97), .IN5(
        product_shift[5]), .IN6(n18), .Q(product2[5]) );
  AO222X1 U18 ( .IN1(N70), .IN2(n100), .IN3(N121), .IN4(n97), .IN5(
        product_shift[49]), .IN6(n18), .Q(product2[50]) );
  AO222X1 U19 ( .IN1(N24), .IN2(n100), .IN3(N75), .IN4(n97), .IN5(
        product_shift[4]), .IN6(n95), .Q(product2[4]) );
  AO222X1 U20 ( .IN1(N69), .IN2(n100), .IN3(N120), .IN4(n97), .IN5(
        product_shift[49]), .IN6(n96), .Q(product2[49]) );
  AO222X1 U21 ( .IN1(N68), .IN2(n100), .IN3(N119), .IN4(n97), .IN5(
        product_shift[48]), .IN6(n18), .Q(product2[48]) );
  AO222X1 U22 ( .IN1(N67), .IN2(n100), .IN3(N118), .IN4(n97), .IN5(
        product_shift[47]), .IN6(n96), .Q(product2[47]) );
  AO222X1 U23 ( .IN1(N66), .IN2(n100), .IN3(N117), .IN4(n97), .IN5(
        product_shift[46]), .IN6(n18), .Q(product2[46]) );
  AO222X1 U24 ( .IN1(N65), .IN2(n100), .IN3(N116), .IN4(n97), .IN5(
        product_shift[45]), .IN6(n95), .Q(product2[45]) );
  AO222X1 U25 ( .IN1(N64), .IN2(n101), .IN3(N115), .IN4(n98), .IN5(
        product_shift[44]), .IN6(n96), .Q(product2[44]) );
  AO222X1 U26 ( .IN1(N63), .IN2(n101), .IN3(N114), .IN4(n98), .IN5(
        product_shift[43]), .IN6(n96), .Q(product2[43]) );
  AO222X1 U27 ( .IN1(N62), .IN2(n101), .IN3(N113), .IN4(n98), .IN5(
        product_shift[42]), .IN6(n96), .Q(product2[42]) );
  AO222X1 U28 ( .IN1(N61), .IN2(n101), .IN3(N112), .IN4(n98), .IN5(
        product_shift[41]), .IN6(n96), .Q(product2[41]) );
  AO222X1 U29 ( .IN1(N60), .IN2(n101), .IN3(N111), .IN4(n98), .IN5(
        product_shift[40]), .IN6(n96), .Q(product2[40]) );
  AO222X1 U30 ( .IN1(N23), .IN2(n101), .IN3(N74), .IN4(n98), .IN5(
        product_shift[3]), .IN6(n96), .Q(product2[3]) );
  AO222X1 U31 ( .IN1(N59), .IN2(n101), .IN3(N110), .IN4(n98), .IN5(
        product_shift[39]), .IN6(n96), .Q(product2[39]) );
  AO222X1 U32 ( .IN1(N58), .IN2(n101), .IN3(N109), .IN4(n98), .IN5(
        product_shift[38]), .IN6(n96), .Q(product2[38]) );
  AO222X1 U33 ( .IN1(N57), .IN2(n101), .IN3(N108), .IN4(n98), .IN5(
        product_shift[37]), .IN6(n96), .Q(product2[37]) );
  AO222X1 U34 ( .IN1(N56), .IN2(n101), .IN3(N107), .IN4(n98), .IN5(
        product_shift[36]), .IN6(n96), .Q(product2[36]) );
  AO222X1 U35 ( .IN1(N55), .IN2(n101), .IN3(N106), .IN4(n98), .IN5(n7), .IN6(
        n96), .Q(product2[35]) );
  AO222X1 U36 ( .IN1(N54), .IN2(n101), .IN3(N105), .IN4(n98), .IN5(n13), .IN6(
        n96), .Q(product2[34]) );
  AO222X1 U37 ( .IN1(N53), .IN2(n102), .IN3(N104), .IN4(n17), .IN5(n26), .IN6(
        n96), .Q(product2[33]) );
  AO222X1 U38 ( .IN1(N52), .IN2(n102), .IN3(N103), .IN4(n17), .IN5(n34), .IN6(
        n18), .Q(product2[32]) );
  AO222X1 U39 ( .IN1(N51), .IN2(n102), .IN3(N102), .IN4(n17), .IN5(n42), .IN6(
        n18), .Q(product2[31]) );
  AO222X1 U40 ( .IN1(N50), .IN2(n102), .IN3(N101), .IN4(n17), .IN5(n48), .IN6(
        n18), .Q(product2[30]) );
  AO222X1 U41 ( .IN1(N22), .IN2(n102), .IN3(N73), .IN4(n17), .IN5(
        product_shift[2]), .IN6(n18), .Q(product2[2]) );
  AO222X1 U42 ( .IN1(N49), .IN2(n102), .IN3(N100), .IN4(n17), .IN5(n55), .IN6(
        n18), .Q(product2[29]) );
  AO222X1 U43 ( .IN1(N48), .IN2(n102), .IN3(N99), .IN4(n17), .IN5(n64), .IN6(
        n18), .Q(product2[28]) );
  AO222X1 U44 ( .IN1(N47), .IN2(n102), .IN3(N98), .IN4(n17), .IN5(n75), .IN6(
        n18), .Q(product2[27]) );
  AO222X1 U45 ( .IN1(N46), .IN2(n102), .IN3(N97), .IN4(n17), .IN5(n86), .IN6(
        n18), .Q(product2[26]) );
  AO222X1 U46 ( .IN1(N45), .IN2(n102), .IN3(N96), .IN4(n17), .IN5(
        product_shift[25]), .IN6(n18), .Q(product2[25]) );
  AO222X1 U48 ( .IN1(N43), .IN2(n102), .IN3(N94), .IN4(n97), .IN5(
        product_shift[23]), .IN6(n18), .Q(product2[23]) );
  AO222X1 U49 ( .IN1(N42), .IN2(n103), .IN3(N93), .IN4(n99), .IN5(
        product_shift[22]), .IN6(n18), .Q(product2[22]) );
  AO222X1 U50 ( .IN1(N41), .IN2(n103), .IN3(N92), .IN4(n99), .IN5(
        product_shift[21]), .IN6(n95), .Q(product2[21]) );
  AO222X1 U51 ( .IN1(N40), .IN2(n103), .IN3(N91), .IN4(n99), .IN5(
        product_shift[20]), .IN6(n95), .Q(product2[20]) );
  AO222X1 U52 ( .IN1(N21), .IN2(n103), .IN3(N72), .IN4(n99), .IN5(n95), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U53 ( .IN1(N39), .IN2(n103), .IN3(N90), .IN4(n99), .IN5(
        product_shift[19]), .IN6(n95), .Q(product2[19]) );
  AO222X1 U54 ( .IN1(N38), .IN2(n103), .IN3(N89), .IN4(n99), .IN5(
        product_shift[18]), .IN6(n95), .Q(product2[18]) );
  AO222X1 U55 ( .IN1(N37), .IN2(n103), .IN3(N88), .IN4(n99), .IN5(
        product_shift[17]), .IN6(n95), .Q(product2[17]) );
  AO222X1 U56 ( .IN1(N36), .IN2(n103), .IN3(N87), .IN4(n99), .IN5(
        product_shift[16]), .IN6(n95), .Q(product2[16]) );
  AO222X1 U57 ( .IN1(N35), .IN2(n103), .IN3(N86), .IN4(n99), .IN5(
        product_shift[15]), .IN6(n95), .Q(product2[15]) );
  AO222X1 U58 ( .IN1(N34), .IN2(n103), .IN3(N85), .IN4(n99), .IN5(
        product_shift[14]), .IN6(n95), .Q(product2[14]) );
  AO222X1 U59 ( .IN1(N33), .IN2(n103), .IN3(N84), .IN4(n99), .IN5(
        product_shift[13]), .IN6(n95), .Q(product2[13]) );
  AO222X1 U60 ( .IN1(N32), .IN2(n103), .IN3(N83), .IN4(n99), .IN5(
        product_shift[12]), .IN6(n95), .Q(product2[12]) );
  AO222X1 U61 ( .IN1(N31), .IN2(n104), .IN3(N82), .IN4(n99), .IN5(
        product_shift[11]), .IN6(n95), .Q(product2[11]) );
  AO222X1 U62 ( .IN1(N30), .IN2(n104), .IN3(N81), .IN4(n98), .IN5(
        product_shift[10]), .IN6(n96), .Q(product2[10]) );
  XOR2X1 U64 ( .IN1(n165), .IN2(product_shift[1]), .Q(n18) );
  AND2X1 U65 ( .IN1(product_shift[1]), .IN2(n165), .Q(n17) );
  AO222X1 U66 ( .IN1(N215), .IN2(n93), .IN3(N138), .IN4(n9), .IN5(N188), .IN6(
        n8), .Q(add_sum[9]) );
  AO222X1 U67 ( .IN1(N214), .IN2(n93), .IN3(N137), .IN4(n9), .IN5(N187), .IN6(
        n8), .Q(add_sum[8]) );
  AO222X1 U68 ( .IN1(N213), .IN2(n93), .IN3(N136), .IN4(n9), .IN5(N186), .IN6(
        n8), .Q(add_sum[7]) );
  AO222X1 U69 ( .IN1(N212), .IN2(n93), .IN3(N135), .IN4(n9), .IN5(N185), .IN6(
        n8), .Q(add_sum[6]) );
  AO222X1 U70 ( .IN1(N211), .IN2(n93), .IN3(N134), .IN4(n9), .IN5(N184), .IN6(
        n8), .Q(add_sum[5]) );
  AO222X1 U71 ( .IN1(N210), .IN2(n93), .IN3(N133), .IN4(n9), .IN5(N183), .IN6(
        n8), .Q(add_sum[4]) );
  AO222X1 U72 ( .IN1(N209), .IN2(n93), .IN3(N132), .IN4(n9), .IN5(N182), .IN6(
        n8), .Q(add_sum[3]) );
  AO222X1 U73 ( .IN1(N208), .IN2(n93), .IN3(N131), .IN4(n9), .IN5(N181), .IN6(
        n8), .Q(add_sum[2]) );
  AO222X1 U74 ( .IN1(N230), .IN2(n93), .IN3(n9), .IN4(N153), .IN5(n8), .IN6(
        N203), .Q(add_sum[24]) );
  AO222X1 U75 ( .IN1(N229), .IN2(n93), .IN3(N152), .IN4(n9), .IN5(n8), .IN6(
        N202), .Q(add_sum[23]) );
  AO222X1 U76 ( .IN1(N228), .IN2(n93), .IN3(N151), .IN4(n9), .IN5(N201), .IN6(
        n8), .Q(add_sum[22]) );
  AO222X1 U77 ( .IN1(N227), .IN2(n93), .IN3(N150), .IN4(n9), .IN5(N200), .IN6(
        n8), .Q(add_sum[21]) );
  AO222X1 U78 ( .IN1(N226), .IN2(n94), .IN3(N149), .IN4(n9), .IN5(N199), .IN6(
        n8), .Q(add_sum[20]) );
  AO222X1 U79 ( .IN1(N207), .IN2(n94), .IN3(N130), .IN4(n9), .IN5(N180), .IN6(
        n8), .Q(add_sum[1]) );
  AO222X1 U80 ( .IN1(N225), .IN2(n94), .IN3(N148), .IN4(n9), .IN5(N198), .IN6(
        n8), .Q(add_sum[19]) );
  AO222X1 U81 ( .IN1(N224), .IN2(n94), .IN3(N147), .IN4(n9), .IN5(N197), .IN6(
        n8), .Q(add_sum[18]) );
  AO222X1 U82 ( .IN1(N223), .IN2(n94), .IN3(N146), .IN4(n9), .IN5(N196), .IN6(
        n8), .Q(add_sum[17]) );
  AO222X1 U83 ( .IN1(N222), .IN2(n94), .IN3(N145), .IN4(n9), .IN5(N195), .IN6(
        n8), .Q(add_sum[16]) );
  AO222X1 U84 ( .IN1(N221), .IN2(n94), .IN3(N144), .IN4(n9), .IN5(N194), .IN6(
        n8), .Q(add_sum[15]) );
  AO222X1 U85 ( .IN1(N220), .IN2(n94), .IN3(N143), .IN4(n9), .IN5(N193), .IN6(
        n8), .Q(add_sum[14]) );
  AO222X1 U86 ( .IN1(N219), .IN2(n94), .IN3(N142), .IN4(n9), .IN5(N192), .IN6(
        n8), .Q(add_sum[13]) );
  AO222X1 U87 ( .IN1(N218), .IN2(n94), .IN3(N141), .IN4(n9), .IN5(N191), .IN6(
        n8), .Q(add_sum[12]) );
  AO222X1 U88 ( .IN1(N217), .IN2(n94), .IN3(N140), .IN4(n9), .IN5(N190), .IN6(
        n8), .Q(add_sum[11]) );
  AO222X1 U89 ( .IN1(N216), .IN2(n94), .IN3(N139), .IN4(n9), .IN5(N189), .IN6(
        n8), .Q(add_sum[10]) );
  AO222X1 U90 ( .IN1(N206), .IN2(n94), .IN3(N129), .IN4(n9), .IN5(N179), .IN6(
        n8), .Q(add_sum[0]) );
  XOR2X1 U92 ( .IN1(add_sign_b), .IN2(add_sign_a), .Q(n22) );
  AO22X1 U94 ( .IN1(add_greater_flag2), .IN2(add_sign_a), .IN3(add_sign_b), 
        .IN4(n166), .Q(add_new_sign) );
  booth2_DW01_sub_0 sub_157 ( .A({1'b0, add_new_b[23:11], n14, n27, n35, n56, 
        n65, n51, n60, n71, n82, n90, n91}), .B({1'b0, add_new_a[23:5], n70, 
        n78, n84, n80, add_new_a[0]}), .CI(1'b0), .DIFF({N230, N229, N228, 
        N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210, N209, N208, N207, N206}) );
  booth2_DW01_sub_1 sub_149 ( .A({1'b0, add_new_a[23:11], n21, n30, n38, n66, 
        n76, n59, n70, n78, n84, n80, n88}), .B({1'b0, add_new_b[23:3], n82, 
        n90, add_new_b[0]}), .CI(1'b0), .DIFF({N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179}) );
  booth2_DW01_add_0 add_96 ( .A({product_shift[49], product_shift[49:36], n7, 
        n13, n26, n34, n42, n48, n55, n64, n75, n86, product_shift[25:0]}), 
        .B({combined_negative_b[24:9], n11, n24, n32, n40, n46, n53, n62, n73, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N121, N120, 
        N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, 
        N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, 
        SYNOPSYS_UNCONNECTED__0, N94, N93, N92, N91, N90, N89, N88, N87, N86, 
        N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth2_DW01_add_1 add_89 ( .A({product_shift[49], product_shift[49:35], n13, 
        n26, n34, n42, n48, n55, n64, n75, n86, product_shift[25:0]}), .B({
        1'b0, combined_b[23:8], n20, n29, n37, n44, n50, n58, n68, 
        combined_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, SYNOPSYS_UNCONNECTED__2, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, SYNOPSYS_UNCONNECTED__3}) );
  booth2_DW01_add_2 r71 ( .A({1'b0, add_new_a[23:11], n21, n30, n38, n66, n76, 
        n59, n70, n78, n84, n80, n88}), .B({1'b0, add_new_b[23:11], n14, n27, 
        n35, n56, n65, n51, n60, n71, n82, n90, n91}), .CI(1'b0), .SUM({N153, 
        N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129}) );
  INVX0 U4 ( .INP(n79), .ZN(n80) );
  NBUFFX2 U5 ( .INP(product_shift[35]), .Z(n7) );
  AO221X1 U8 ( .IN1(n21), .IN2(n150), .IN3(add_new_a[11]), .IN4(n151), .IN5(
        n128), .Q(n129) );
  AND2X2 U12 ( .IN1(N124), .IN2(n22), .Q(n8) );
  XNOR2X1 U47 ( .IN1(add_sign_a), .IN2(add_sign_b), .Q(n9) );
  OA221X1 U63 ( .IN1(add_new_a[12]), .IN2(n152), .IN3(add_new_a[11]), .IN4(
        n151), .IN5(n129), .Q(n130) );
  INVX0 U91 ( .INP(combined_negative_b[8]), .ZN(n10) );
  INVX0 U93 ( .INP(n10), .ZN(n11) );
  INVX0 U95 ( .INP(product_shift[34]), .ZN(n12) );
  INVX0 U96 ( .INP(n12), .ZN(n13) );
  INVX0 U97 ( .INP(n150), .ZN(n14) );
  INVX0 U98 ( .INP(combined_b[7]), .ZN(n15) );
  INVX0 U99 ( .INP(n15), .ZN(n20) );
  NBUFFX2 U100 ( .INP(add_new_a[10]), .Z(n21) );
  INVX0 U101 ( .INP(combined_negative_b[7]), .ZN(n23) );
  INVX0 U102 ( .INP(n23), .ZN(n24) );
  INVX0 U103 ( .INP(product_shift[33]), .ZN(n25) );
  INVX0 U104 ( .INP(n25), .ZN(n26) );
  INVX0 U105 ( .INP(n149), .ZN(n27) );
  INVX0 U106 ( .INP(combined_b[6]), .ZN(n28) );
  INVX0 U107 ( .INP(n28), .ZN(n29) );
  NBUFFX2 U108 ( .INP(add_new_a[9]), .Z(n30) );
  INVX0 U109 ( .INP(combined_negative_b[6]), .ZN(n31) );
  INVX0 U110 ( .INP(n31), .ZN(n32) );
  INVX0 U111 ( .INP(product_shift[32]), .ZN(n33) );
  INVX0 U112 ( .INP(n33), .ZN(n34) );
  INVX0 U113 ( .INP(n148), .ZN(n35) );
  INVX0 U114 ( .INP(combined_b[5]), .ZN(n36) );
  INVX0 U115 ( .INP(n36), .ZN(n37) );
  NBUFFX2 U116 ( .INP(add_new_a[8]), .Z(n38) );
  INVX0 U117 ( .INP(combined_negative_b[5]), .ZN(n39) );
  INVX0 U118 ( .INP(n39), .ZN(n40) );
  INVX0 U119 ( .INP(product_shift[31]), .ZN(n41) );
  INVX0 U120 ( .INP(n41), .ZN(n42) );
  INVX0 U121 ( .INP(combined_b[4]), .ZN(n43) );
  INVX0 U122 ( .INP(n43), .ZN(n44) );
  INVX0 U123 ( .INP(combined_negative_b[4]), .ZN(n45) );
  INVX0 U124 ( .INP(n45), .ZN(n46) );
  INVX0 U125 ( .INP(product_shift[30]), .ZN(n47) );
  INVX0 U126 ( .INP(n47), .ZN(n48) );
  INVX0 U127 ( .INP(combined_b[3]), .ZN(n49) );
  INVX0 U128 ( .INP(n49), .ZN(n50) );
  INVX0 U129 ( .INP(n145), .ZN(n51) );
  INVX0 U130 ( .INP(combined_negative_b[3]), .ZN(n52) );
  INVX0 U131 ( .INP(n52), .ZN(n53) );
  INVX0 U132 ( .INP(product_shift[29]), .ZN(n54) );
  INVX0 U133 ( .INP(n54), .ZN(n55) );
  INVX0 U134 ( .INP(n147), .ZN(n56) );
  INVX0 U135 ( .INP(combined_b[2]), .ZN(n57) );
  INVX0 U136 ( .INP(n57), .ZN(n58) );
  NBUFFX2 U137 ( .INP(add_new_a[5]), .Z(n59) );
  INVX0 U138 ( .INP(n144), .ZN(n60) );
  INVX0 U139 ( .INP(combined_negative_b[2]), .ZN(n61) );
  INVX0 U140 ( .INP(n61), .ZN(n62) );
  INVX0 U141 ( .INP(product_shift[28]), .ZN(n63) );
  INVX0 U142 ( .INP(n63), .ZN(n64) );
  INVX0 U143 ( .INP(n146), .ZN(n65) );
  NBUFFX2 U144 ( .INP(add_new_a[7]), .Z(n66) );
  INVX0 U145 ( .INP(combined_b[1]), .ZN(n67) );
  INVX0 U146 ( .INP(n67), .ZN(n68) );
  INVX0 U147 ( .INP(add_new_a[4]), .ZN(n69) );
  INVX0 U148 ( .INP(n69), .ZN(n70) );
  INVX0 U149 ( .INP(n143), .ZN(n71) );
  INVX0 U150 ( .INP(combined_negative_b[1]), .ZN(n72) );
  INVX0 U151 ( .INP(n72), .ZN(n73) );
  INVX0 U152 ( .INP(product_shift[27]), .ZN(n74) );
  INVX0 U153 ( .INP(n74), .ZN(n75) );
  NBUFFX2 U154 ( .INP(add_new_a[6]), .Z(n76) );
  INVX0 U155 ( .INP(add_new_a[3]), .ZN(n77) );
  INVX0 U156 ( .INP(n77), .ZN(n78) );
  DELLN1X2 U157 ( .INP(add_new_b[0]), .Z(n91) );
  NBUFFX2 U158 ( .INP(n19), .Z(n94) );
  NBUFFX2 U159 ( .INP(n19), .Z(n93) );
  NBUFFX2 U160 ( .INP(n92), .Z(n105) );
  NBUFFX2 U161 ( .INP(n92), .Z(n106) );
  NBUFFX2 U162 ( .INP(n92), .Z(n107) );
  NBUFFX2 U163 ( .INP(n92), .Z(n108) );
  NBUFFX2 U164 ( .INP(n92), .Z(n109) );
  NBUFFX2 U165 ( .INP(n92), .Z(n110) );
  NBUFFX2 U166 ( .INP(n92), .Z(n111) );
  NBUFFX2 U167 ( .INP(n92), .Z(n112) );
  NBUFFX2 U168 ( .INP(n92), .Z(n113) );
  NBUFFX2 U169 ( .INP(n92), .Z(n115) );
  NBUFFX2 U170 ( .INP(n92), .Z(n116) );
  NBUFFX2 U171 ( .INP(n92), .Z(n114) );
  NBUFFX2 U172 ( .INP(n92), .Z(n117) );
  NOR2X0 U173 ( .IN1(n9), .IN2(n8), .QN(n19) );
  INVX0 U174 ( .INP(n88), .ZN(n164) );
  NBUFFX2 U175 ( .INP(n16), .Z(n103) );
  NBUFFX2 U176 ( .INP(n16), .Z(n101) );
  NBUFFX2 U177 ( .INP(n16), .Z(n100) );
  NBUFFX2 U178 ( .INP(n16), .Z(n102) );
  NBUFFX2 U179 ( .INP(n16), .Z(n104) );
  NBUFFX2 U180 ( .INP(n18), .Z(n95) );
  NBUFFX2 U181 ( .INP(n18), .Z(n96) );
  NBUFFX2 U182 ( .INP(n17), .Z(n99) );
  NBUFFX2 U183 ( .INP(n17), .Z(n98) );
  NBUFFX2 U184 ( .INP(n17), .Z(n97) );
  NBUFFX2 U185 ( .INP(reset), .Z(n92) );
  INVX0 U186 ( .INP(n87), .ZN(n88) );
  OA222X1 U187 ( .IN1(n84), .IN2(n81), .IN3(n80), .IN4(n119), .IN5(n118), 
        .IN6(n89), .Q(n120) );
  INVX0 U188 ( .INP(add_new_b[3]), .ZN(n143) );
  INVX0 U189 ( .INP(add_new_b[8]), .ZN(n148) );
  INVX0 U190 ( .INP(add_new_b[14]), .ZN(n154) );
  INVX0 U191 ( .INP(add_new_b[20]), .ZN(n160) );
  INVX0 U192 ( .INP(add_new_b[5]), .ZN(n145) );
  INVX0 U193 ( .INP(add_new_b[11]), .ZN(n151) );
  INVX0 U194 ( .INP(add_new_b[17]), .ZN(n157) );
  INVX0 U195 ( .INP(add_new_b[22]), .ZN(n162) );
  INVX0 U196 ( .INP(add_new_b[7]), .ZN(n147) );
  INVX0 U197 ( .INP(add_new_b[9]), .ZN(n149) );
  INVX0 U198 ( .INP(add_new_b[10]), .ZN(n150) );
  INVX0 U199 ( .INP(add_new_b[4]), .ZN(n144) );
  INVX0 U200 ( .INP(add_new_b[6]), .ZN(n146) );
  INVX0 U201 ( .INP(add_new_b[12]), .ZN(n152) );
  NOR2X0 U202 ( .IN1(n165), .IN2(product_shift[1]), .QN(n16) );
  INVX0 U203 ( .INP(add_new_b[13]), .ZN(n153) );
  INVX0 U204 ( .INP(add_new_b[15]), .ZN(n155) );
  INVX0 U205 ( .INP(add_new_b[19]), .ZN(n159) );
  INVX0 U206 ( .INP(add_new_b[21]), .ZN(n161) );
  INVX0 U207 ( .INP(add_new_b[16]), .ZN(n156) );
  INVX0 U208 ( .INP(add_new_b[18]), .ZN(n158) );
  INVX0 U209 ( .INP(add_new_b[23]), .ZN(n163) );
  INVX0 U210 ( .INP(product_shift[0]), .ZN(n165) );
  INVX0 U211 ( .INP(add_greater_flag2), .ZN(n166) );
  INVX0 U213 ( .INP(add_new_a[1]), .ZN(n79) );
  INVX0 U214 ( .INP(add_new_b[2]), .ZN(n81) );
  INVX0 U215 ( .INP(n81), .ZN(n82) );
  INVX0 U216 ( .INP(add_new_a[2]), .ZN(n83) );
  INVX0 U217 ( .INP(n83), .ZN(n84) );
  INVX0 U218 ( .INP(product_shift[26]), .ZN(n85) );
  INVX0 U219 ( .INP(n85), .ZN(n86) );
  INVX0 U220 ( .INP(add_new_a[0]), .ZN(n87) );
  INVX0 U221 ( .INP(add_new_b[1]), .ZN(n89) );
  INVX0 U222 ( .INP(n89), .ZN(n90) );
  AND2X1 U223 ( .IN1(n162), .IN2(add_new_a[22]), .Q(n141) );
  NOR2X0 U224 ( .IN1(n164), .IN2(n91), .QN(n118) );
  AND2X1 U225 ( .IN1(n89), .IN2(n118), .Q(n119) );
  AO221X1 U226 ( .IN1(n84), .IN2(n81), .IN3(n78), .IN4(n143), .IN5(n120), .Q(
        n121) );
  OA221X1 U227 ( .IN1(n70), .IN2(n144), .IN3(n78), .IN4(n143), .IN5(n121), .Q(
        n122) );
  AO221X1 U228 ( .IN1(n70), .IN2(n144), .IN3(n59), .IN4(n145), .IN5(n122), .Q(
        n123) );
  OA221X1 U229 ( .IN1(n76), .IN2(n146), .IN3(n59), .IN4(n145), .IN5(n123), .Q(
        n124) );
  AO221X1 U230 ( .IN1(n76), .IN2(n146), .IN3(n66), .IN4(n147), .IN5(n124), .Q(
        n125) );
  OA221X1 U231 ( .IN1(n38), .IN2(n148), .IN3(n66), .IN4(n147), .IN5(n125), .Q(
        n126) );
  AO221X1 U232 ( .IN1(n38), .IN2(n148), .IN3(n30), .IN4(n149), .IN5(n126), .Q(
        n127) );
  OA221X1 U233 ( .IN1(n30), .IN2(n149), .IN3(n21), .IN4(n150), .IN5(n127), .Q(
        n128) );
  AO221X1 U234 ( .IN1(add_new_a[12]), .IN2(n152), .IN3(add_new_a[13]), .IN4(
        n153), .IN5(n130), .Q(n131) );
  OA221X1 U235 ( .IN1(add_new_a[14]), .IN2(n154), .IN3(add_new_a[13]), .IN4(
        n153), .IN5(n131), .Q(n132) );
  AO221X1 U236 ( .IN1(add_new_a[14]), .IN2(n154), .IN3(add_new_a[15]), .IN4(
        n155), .IN5(n132), .Q(n133) );
  OA221X1 U237 ( .IN1(add_new_a[16]), .IN2(n156), .IN3(add_new_a[15]), .IN4(
        n155), .IN5(n133), .Q(n134) );
  AO221X1 U238 ( .IN1(add_new_a[16]), .IN2(n156), .IN3(add_new_a[17]), .IN4(
        n157), .IN5(n134), .Q(n135) );
  OA221X1 U239 ( .IN1(add_new_a[18]), .IN2(n158), .IN3(add_new_a[17]), .IN4(
        n157), .IN5(n135), .Q(n136) );
  AO221X1 U240 ( .IN1(add_new_a[18]), .IN2(n158), .IN3(add_new_a[19]), .IN4(
        n159), .IN5(n136), .Q(n137) );
  OA221X1 U241 ( .IN1(add_new_a[20]), .IN2(n160), .IN3(add_new_a[19]), .IN4(
        n159), .IN5(n137), .Q(n138) );
  AO221X1 U242 ( .IN1(add_new_a[20]), .IN2(n160), .IN3(add_new_a[21]), .IN4(
        n161), .IN5(n138), .Q(n139) );
  OA221X1 U243 ( .IN1(add_new_a[22]), .IN2(n162), .IN3(add_new_a[21]), .IN4(
        n161), .IN5(n139), .Q(n140) );
  OA22X1 U244 ( .IN1(add_new_a[23]), .IN2(n163), .IN3(n141), .IN4(n140), .Q(
        n142) );
  AO21X1 U245 ( .IN1(add_new_a[23]), .IN2(n163), .IN3(n142), .Q(N124) );
endmodule


module booth3_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(SUM[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module booth3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n22), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  NAND2X0 U1 ( .IN1(A[49]), .IN2(carry[49]), .QN(n1) );
  XOR3X1 U2 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U3 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U4 ( .IN1(B[49]), .IN2(carry[49]), .QN(n2) );
  NAND2X1 U5 ( .IN1(B[49]), .IN2(A[49]), .QN(n3) );
  NAND3X0 U6 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[50]) );
  XOR3X1 U7 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U8 ( .IN1(A[46]), .IN2(carry[46]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[46]), .IN2(carry[46]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[46]), .IN2(A[46]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[47]) );
  DELLN2X2 U12 ( .INP(carry[45]), .Z(n7) );
  XOR3X2 U13 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U14 ( .IN1(A[44]), .IN2(B[44]), .QN(n8) );
  NAND2X0 U15 ( .IN1(A[44]), .IN2(carry[44]), .QN(n9) );
  NAND2X0 U16 ( .IN1(B[44]), .IN2(carry[44]), .QN(n10) );
  NAND3X0 U17 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[45]) );
  XOR2X1 U18 ( .IN1(A[45]), .IN2(B[45]), .Q(n11) );
  XOR2X1 U19 ( .IN1(n11), .IN2(n7), .Q(SUM[45]) );
  NAND2X0 U20 ( .IN1(A[45]), .IN2(B[45]), .QN(n12) );
  NAND2X0 U21 ( .IN1(A[45]), .IN2(carry[45]), .QN(n13) );
  NAND2X0 U22 ( .IN1(B[45]), .IN2(carry[45]), .QN(n14) );
  NAND3X0 U23 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U24 ( .IN1(A[47]), .IN2(B[47]), .QN(n15) );
  NAND2X0 U25 ( .IN1(A[47]), .IN2(carry[47]), .QN(n16) );
  NAND2X0 U26 ( .IN1(B[47]), .IN2(carry[47]), .QN(n17) );
  NAND3X0 U27 ( .IN1(n16), .IN2(n17), .IN3(n15), .QN(carry[48]) );
  XOR2X1 U28 ( .IN1(A[48]), .IN2(B[48]), .Q(n18) );
  XOR2X1 U29 ( .IN1(n18), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U30 ( .IN1(A[48]), .IN2(B[48]), .QN(n19) );
  NAND2X0 U31 ( .IN1(A[48]), .IN2(carry[48]), .QN(n20) );
  NAND2X0 U32 ( .IN1(B[48]), .IN2(carry[48]), .QN(n21) );
  NAND3X0 U33 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[49]) );
  AND2X1 U34 ( .IN1(A[26]), .IN2(B[26]), .Q(n22) );
  XOR2X1 U35 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n22), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X1 U2 ( .IN1(A[43]), .IN2(B[43]), .QN(n1) );
  NAND2X1 U3 ( .IN1(A[43]), .IN2(carry[43]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[43]), .IN2(carry[43]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[44]) );
  XOR2X1 U6 ( .IN1(A[44]), .IN2(B[44]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[44]), .Q(SUM[44]) );
  NAND2X0 U8 ( .IN1(A[44]), .IN2(B[44]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[44]), .IN2(carry[44]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[44]), .IN2(carry[44]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[45]) );
  XOR3X2 U12 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(B[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[48]), .IN2(carry[48]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[48]), .IN2(carry[48]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[49]) );
  XOR2X1 U17 ( .IN1(A[49]), .IN2(B[49]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(B[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[49]), .IN2(carry[49]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[49]), .IN2(carry[49]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[50]) );
  XOR3X2 U23 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U24 ( .IN1(A[46]), .IN2(B[46]), .QN(n15) );
  NAND2X0 U25 ( .IN1(A[46]), .IN2(carry[46]), .QN(n16) );
  NAND2X0 U26 ( .IN1(B[46]), .IN2(carry[46]), .QN(n17) );
  NAND3X0 U27 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[47]) );
  XOR2X1 U28 ( .IN1(A[47]), .IN2(B[47]), .Q(n18) );
  XOR2X1 U29 ( .IN1(n18), .IN2(carry[47]), .Q(SUM[47]) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U32 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U33 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[48]) );
  AND2X1 U34 ( .IN1(A[26]), .IN2(B[26]), .Q(n22) );
  XOR2X1 U35 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth3_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[7]), .IN2(A[7]), .Q(SUM[7]) );
endmodule


module booth3 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_sign_a, add_sign_b, add_sum, 
        add_new_exponent, add_updated_exponent_o, add_updated_add_sum_o, 
        add_exception1_o, add_exception2_o, add_new_sign, add_new_sign2, 
        add_sign_a5, add_sign_b5, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [24:0] add_sum;
  input [7:0] add_new_exponent;
  output [7:0] add_updated_exponent_o;
  output [24:0] add_updated_add_sum_o;
  input clk, reset, new_sign, add_sign_a, add_sign_b, add_new_sign, s;
  output new_sign2, add_exception1_o, add_exception2_o, add_new_sign2,
         add_sign_a5, add_sign_b5, s2;
  wire   N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146,
         N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, add_exception1, add_exception2, N192,
         N193, N194, N195, N196, N197, N198, N199, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N298,
         N299, N300, N301, N302, N303, N304, N340, N342, N343, N344, N345,
         N346, N347, N383, N384, N385, N386, N387, N388, N389, N424, N426,
         N427, N428, N429, N430, N464, N465, N466, N467, N468, N469, N470,
         N504, N505, N506, N507, N508, N509, N541, N542, N543, N544, N545,
         N546, N547, N580, N582, N583, N584, N585, N615, N616, N617, N618,
         N619, N620, N621, N651, N652, N653, N654, N655, N656, N684, N685,
         N686, N687, N688, N689, N690, N719, N720, N721, N722, N723, N749,
         N750, N751, N752, N753, N754, N755, N781, N782, N783, N784, N785,
         N786, N810, N811, N812, N813, N814, N815, N816, N841, N843, N844,
         N845, N867, N868, N869, N870, N871, N872, N873, N895, N896, N897,
         N898, N899, N900, N920, N921, N922, N923, N924, N925, N926, N947,
         N948, N949, N950, N951, N969, N970, N971, N972, N973, N974, N975,
         N993, N994, N995, N996, N997, N998, N1014, N1015, N1016, N1017, N1018,
         N1019, N1020, \sub_595/carry[2] , \sub_595/carry[3] ,
         \sub_595/carry[4] , \sub_595/carry[5] , \sub_595/carry[6] ,
         \sub_595/carry[7] , \sub_579/carry[7] , \sub_579/carry[6] ,
         \sub_579/carry[5] , \sub_579/carry[4] , \sub_579/carry[3] ,
         \sub_563/carry[2] , \sub_563/carry[3] , \sub_563/carry[4] ,
         \sub_563/carry[5] , \sub_563/carry[6] , \sub_563/carry[7] ,
         \sub_547/carry[7] , \sub_547/carry[6] , \sub_547/carry[5] ,
         \sub_547/carry[4] , \sub_531/carry[2] , \sub_531/carry[3] ,
         \sub_531/carry[4] , \sub_531/carry[5] , \sub_531/carry[6] ,
         \sub_531/carry[7] , \sub_515/carry[7] , \sub_515/carry[6] ,
         \sub_515/carry[5] , \sub_515/carry[4] , \sub_515/carry[3] ,
         \sub_499/carry[2] , \sub_499/carry[3] , \sub_499/carry[4] ,
         \sub_499/carry[5] , \sub_499/carry[6] , \sub_499/carry[7] ,
         \sub_483/carry[7] , \sub_483/carry[6] , \sub_467/carry[2] ,
         \sub_467/carry[3] , \sub_467/carry[4] , \sub_467/carry[5] ,
         \sub_467/carry[6] , \sub_467/carry[7] , \sub_451/carry[7] ,
         \sub_451/carry[6] , \sub_451/carry[5] , \sub_451/carry[4] ,
         \sub_451/carry[3] , \sub_435/carry[2] , \sub_435/carry[3] ,
         \sub_435/carry[4] , \sub_435/carry[5] , \sub_435/carry[6] ,
         \sub_435/carry[7] , \sub_419/carry[7] , \sub_419/carry[6] ,
         \sub_419/carry[5] , \sub_419/carry[4] , \sub_403/carry[2] ,
         \sub_403/carry[3] , \sub_403/carry[4] , \sub_403/carry[5] ,
         \sub_403/carry[6] , \sub_403/carry[7] , \sub_387/carry[7] ,
         \sub_387/carry[6] , \sub_387/carry[5] , \sub_387/carry[4] ,
         \sub_387/carry[3] , \sub_371/carry[2] , \sub_371/carry[3] ,
         \sub_371/carry[4] , \sub_371/carry[5] , \sub_371/carry[6] ,
         \sub_371/carry[7] , \sub_355/carry[7] , \sub_355/carry[6] ,
         \sub_355/carry[5] , \sub_339/carry[2] , \sub_339/carry[3] ,
         \sub_339/carry[4] , \sub_339/carry[5] , \sub_339/carry[6] ,
         \sub_339/carry[7] , \sub_323/carry[7] , \sub_323/carry[6] ,
         \sub_323/carry[5] , \sub_323/carry[4] , \sub_323/carry[3] ,
         \sub_307/carry[2] , \sub_307/carry[3] , \sub_307/carry[4] ,
         \sub_307/carry[5] , \sub_307/carry[6] , \sub_307/carry[7] ,
         \sub_291/carry[7] , \sub_291/carry[6] , \sub_291/carry[5] ,
         \sub_291/carry[4] , \sub_275/carry[2] , \sub_275/carry[3] ,
         \sub_275/carry[4] , \sub_275/carry[5] , \sub_275/carry[6] ,
         \sub_275/carry[7] , \sub_259/carry[7] , \sub_259/carry[6] ,
         \sub_259/carry[5] , \sub_259/carry[4] , \sub_259/carry[3] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   [24:0] add_updated_add_sum;
  wire   [7:0] add_updated_exponent;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[23] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];
  assign N340 = add_new_exponent[0];
  assign N424 = add_new_exponent[1];
  assign N580 = add_new_exponent[2];
  assign N841 = add_new_exponent[3];

  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n100), .Q(new_sign2)
         );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n100), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n100), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n100), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n100), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n99), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n98), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n97), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n96), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n96), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n95), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n94), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n94), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(n4), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n16), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n22), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n28), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n34), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n40), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n47), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n94), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n93), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n92), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n92), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n92), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n92), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n92), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n2), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n8), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n14), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n20), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n26), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n32), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n38), .CLK(clk), .RSTB(n92), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n91), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n91), 
        .Q(new_exponent2[0]) );
  DFFARX1 add_sign_a5_reg ( .D(add_sign_a), .CLK(clk), .RSTB(n91), .Q(
        add_sign_a5) );
  DFFARX1 add_sign_b5_reg ( .D(add_sign_b), .CLK(clk), .RSTB(n91), .Q(
        add_sign_b5) );
  DFFARX1 \add_updated_add_sum_o_reg[24]  ( .D(add_updated_add_sum[24]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[24]) );
  DFFARX1 \add_updated_add_sum_o_reg[23]  ( .D(add_updated_add_sum[23]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[23]) );
  DFFARX1 \add_updated_add_sum_o_reg[22]  ( .D(add_updated_add_sum[22]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[22]) );
  DFFARX1 \add_updated_add_sum_o_reg[21]  ( .D(add_updated_add_sum[21]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[21]) );
  DFFARX1 \add_updated_add_sum_o_reg[20]  ( .D(add_updated_add_sum[20]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[20]) );
  DFFARX1 \add_updated_add_sum_o_reg[19]  ( .D(add_updated_add_sum[19]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[19]) );
  DFFARX1 \add_updated_add_sum_o_reg[18]  ( .D(add_updated_add_sum[18]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[18]) );
  DFFARX1 \add_updated_add_sum_o_reg[17]  ( .D(add_updated_add_sum[17]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[17]) );
  DFFARX1 \add_updated_add_sum_o_reg[16]  ( .D(add_updated_add_sum[16]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[16]) );
  DFFARX1 \add_updated_add_sum_o_reg[15]  ( .D(add_updated_add_sum[15]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[15]) );
  DFFARX1 \add_updated_add_sum_o_reg[14]  ( .D(add_updated_add_sum[14]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[14]) );
  DFFARX1 \add_updated_add_sum_o_reg[13]  ( .D(add_updated_add_sum[13]), .CLK(
        clk), .RSTB(n90), .Q(add_updated_add_sum_o[13]) );
  DFFARX1 \add_updated_add_sum_o_reg[12]  ( .D(add_updated_add_sum[12]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[12]) );
  DFFARX1 \add_updated_add_sum_o_reg[11]  ( .D(add_updated_add_sum[11]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[11]) );
  DFFARX1 \add_updated_add_sum_o_reg[10]  ( .D(add_updated_add_sum[10]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[10]) );
  DFFARX1 \add_updated_add_sum_o_reg[9]  ( .D(add_updated_add_sum[9]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[9]) );
  DFFARX1 \add_updated_add_sum_o_reg[8]  ( .D(add_updated_add_sum[8]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[8]) );
  DFFARX1 \add_updated_add_sum_o_reg[7]  ( .D(add_updated_add_sum[7]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[7]) );
  DFFARX1 \add_updated_add_sum_o_reg[6]  ( .D(add_updated_add_sum[6]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[6]) );
  DFFARX1 \add_updated_add_sum_o_reg[5]  ( .D(add_updated_add_sum[5]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[5]) );
  DFFARX1 \add_updated_add_sum_o_reg[4]  ( .D(add_updated_add_sum[4]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[4]) );
  DFFARX1 \add_updated_add_sum_o_reg[3]  ( .D(add_updated_add_sum[3]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[3]) );
  DFFARX1 \add_updated_add_sum_o_reg[2]  ( .D(add_updated_add_sum[2]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[2]) );
  DFFARX1 \add_updated_add_sum_o_reg[1]  ( .D(add_updated_add_sum[1]), .CLK(
        clk), .RSTB(n89), .Q(add_updated_add_sum_o[1]) );
  DFFARX1 \add_updated_add_sum_o_reg[0]  ( .D(add_updated_add_sum[0]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_add_sum_o[0]) );
  DFFARX1 \add_updated_exponent_o_reg[7]  ( .D(add_updated_exponent[7]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[7]) );
  DFFARX1 \add_updated_exponent_o_reg[6]  ( .D(add_updated_exponent[6]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[6]) );
  DFFARX1 \add_updated_exponent_o_reg[5]  ( .D(add_updated_exponent[5]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[5]) );
  DFFARX1 \add_updated_exponent_o_reg[4]  ( .D(add_updated_exponent[4]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[4]) );
  DFFARX1 \add_updated_exponent_o_reg[3]  ( .D(add_updated_exponent[3]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[3]) );
  DFFARX1 \add_updated_exponent_o_reg[2]  ( .D(add_updated_exponent[2]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[2]) );
  DFFARX1 \add_updated_exponent_o_reg[1]  ( .D(add_updated_exponent[1]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[1]) );
  DFFARX1 \add_updated_exponent_o_reg[0]  ( .D(add_updated_exponent[0]), .CLK(
        clk), .RSTB(n88), .Q(add_updated_exponent_o[0]) );
  DFFARX1 add_exception1_o_reg ( .D(add_exception1), .CLK(clk), .RSTB(n88), 
        .Q(add_exception1_o) );
  DFFARX1 add_exception2_o_reg ( .D(add_exception2), .CLK(clk), .RSTB(n88), 
        .Q(add_exception2_o) );
  DFFARX1 add_new_sign2_reg ( .D(add_new_sign), .CLK(clk), .RSTB(n88), .Q(
        add_new_sign2) );
  booth3_DW01_inc_0 add_203 ( .A({1'b0, add_sum[24:1]}), .SUM({N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201}) );
  booth3_DW01_add_0 add_97 ( .A({product_shift[49], product_shift[49:35], n6, 
        n12, n18, n24, n30, n36, n42, n49, n51, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n2, n8, n14, n20, n26, n32, n38, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N174, N173, 
        N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, 
        N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, 
        N148, SYNOPSYS_UNCONNECTED__0, N146, N145, N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, SYNOPSYS_UNCONNECTED__1}) );
  booth3_DW01_add_1 add_90 ( .A({product_shift[49], product_shift[49:35], n6, 
        n12, n18, n24, n30, n36, n42, n49, n51, product_shift[25:0]}), .B({
        combined_b[24:9], n4, n10, n16, n22, n28, n34, n40, n47, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N123, N122, N121, N120, N119, N118, 
        N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        SYNOPSYS_UNCONNECTED__2, N95, N94, N93, N92, N91, N90, N89, N88, N87, 
        N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        SYNOPSYS_UNCONNECTED__3}) );
  booth3_DW01_inc_1 r235 ( .A({n87, n85, add_new_exponent[5], n78, n75, n71, 
        n68, n65}), .SUM({N199, N198, N197, N196, N195, N194, N193, N192}) );
  XOR2X1 U3 ( .IN1(n74), .IN2(n70), .Q(N781) );
  AO222X1 U4 ( .IN1(N869), .IN2(n129), .IN3(N812), .IN4(n130), .IN5(N841), 
        .IN6(n128), .Q(n190) );
  XNOR2X1 U5 ( .IN1(n77), .IN2(\sub_387/carry[3] ), .Q(N652) );
  XOR2X1 U6 ( .IN1(\sub_419/carry[4] ), .IN2(n81), .Q(N720) );
  XNOR2X1 U7 ( .IN1(n74), .IN2(n77), .Q(N426) );
  XOR2X1 U8 ( .IN1(\sub_467/carry[4] ), .IN2(n81), .Q(N813) );
  NAND2X1 U9 ( .IN1(n70), .IN2(n67), .QN(\sub_371/carry[2] ) );
  XNOR2X1 U10 ( .IN1(n77), .IN2(\sub_451/carry[3] ), .Q(N782) );
  XNOR2X1 U11 ( .IN1(n81), .IN2(\sub_531/carry[4] ), .Q(N923) );
  XOR2X1 U12 ( .IN1(n74), .IN2(n70), .Q(N993) );
  XNOR2X1 U13 ( .IN1(n81), .IN2(\sub_547/carry[4] ), .Q(N948) );
  INVX0 U14 ( .INP(combined_negative_b[7]), .ZN(n1) );
  INVX0 U15 ( .INP(n1), .ZN(n2) );
  INVX0 U16 ( .INP(combined_b[8]), .ZN(n3) );
  INVX0 U17 ( .INP(n3), .ZN(n4) );
  INVX0 U18 ( .INP(product_shift[34]), .ZN(n5) );
  INVX0 U19 ( .INP(n5), .ZN(n6) );
  INVX0 U20 ( .INP(combined_negative_b[6]), .ZN(n7) );
  INVX0 U21 ( .INP(n7), .ZN(n8) );
  INVX0 U22 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U23 ( .INP(n9), .ZN(n10) );
  INVX0 U24 ( .INP(product_shift[33]), .ZN(n11) );
  INVX0 U25 ( .INP(n11), .ZN(n12) );
  INVX0 U26 ( .INP(combined_negative_b[5]), .ZN(n13) );
  INVX0 U27 ( .INP(n13), .ZN(n14) );
  INVX0 U28 ( .INP(combined_b[6]), .ZN(n15) );
  INVX0 U29 ( .INP(n15), .ZN(n16) );
  INVX0 U30 ( .INP(product_shift[32]), .ZN(n17) );
  INVX0 U31 ( .INP(n17), .ZN(n18) );
  INVX0 U32 ( .INP(combined_negative_b[4]), .ZN(n19) );
  INVX0 U33 ( .INP(n19), .ZN(n20) );
  INVX0 U34 ( .INP(combined_b[5]), .ZN(n21) );
  INVX0 U35 ( .INP(n21), .ZN(n22) );
  INVX0 U36 ( .INP(product_shift[31]), .ZN(n23) );
  INVX0 U37 ( .INP(n23), .ZN(n24) );
  INVX0 U38 ( .INP(combined_negative_b[3]), .ZN(n25) );
  INVX0 U39 ( .INP(n25), .ZN(n26) );
  INVX0 U40 ( .INP(combined_b[4]), .ZN(n27) );
  INVX0 U41 ( .INP(n27), .ZN(n28) );
  INVX0 U42 ( .INP(product_shift[30]), .ZN(n29) );
  INVX0 U43 ( .INP(n29), .ZN(n30) );
  INVX0 U44 ( .INP(combined_negative_b[2]), .ZN(n31) );
  INVX0 U45 ( .INP(n31), .ZN(n32) );
  INVX0 U46 ( .INP(combined_b[3]), .ZN(n33) );
  INVX0 U47 ( .INP(n33), .ZN(n34) );
  INVX0 U48 ( .INP(product_shift[29]), .ZN(n35) );
  INVX0 U49 ( .INP(n35), .ZN(n36) );
  INVX0 U50 ( .INP(combined_negative_b[1]), .ZN(n37) );
  INVX0 U51 ( .INP(n37), .ZN(n38) );
  INVX0 U52 ( .INP(combined_b[2]), .ZN(n39) );
  INVX0 U53 ( .INP(n39), .ZN(n40) );
  INVX0 U54 ( .INP(product_shift[28]), .ZN(n41) );
  INVX0 U55 ( .INP(n41), .ZN(n42) );
  INVX0 U56 ( .INP(combined_b[1]), .ZN(n43) );
  INVX0 U57 ( .INP(n43), .ZN(n47) );
  INVX0 U58 ( .INP(product_shift[27]), .ZN(n48) );
  INVX0 U59 ( .INP(n48), .ZN(n49) );
  INVX0 U60 ( .INP(n102), .ZN(n107) );
  INVX0 U61 ( .INP(n104), .ZN(n109) );
  INVX0 U62 ( .INP(n103), .ZN(n108) );
  INVX0 U63 ( .INP(n105), .ZN(n110) );
  NBUFFX2 U64 ( .INP(n116), .Z(n62) );
  NBUFFX2 U65 ( .INP(n233), .Z(n64) );
  NBUFFX2 U66 ( .INP(n52), .Z(n88) );
  NBUFFX2 U67 ( .INP(n52), .Z(n89) );
  NBUFFX2 U68 ( .INP(n52), .Z(n90) );
  NBUFFX2 U69 ( .INP(n52), .Z(n91) );
  NBUFFX2 U70 ( .INP(n52), .Z(n92) );
  NBUFFX2 U71 ( .INP(n52), .Z(n93) );
  NBUFFX2 U72 ( .INP(n52), .Z(n94) );
  NBUFFX2 U73 ( .INP(n52), .Z(n95) );
  NBUFFX2 U77 ( .INP(n52), .Z(n96) );
  NBUFFX2 U78 ( .INP(n52), .Z(n98) );
  NBUFFX2 U79 ( .INP(n52), .Z(n99) );
  NBUFFX2 U80 ( .INP(n52), .Z(n97) );
  NBUFFX2 U81 ( .INP(n52), .Z(n100) );
  INVX0 U82 ( .INP(n67), .ZN(n65) );
  INVX0 U83 ( .INP(n77), .ZN(n76) );
  INVX0 U84 ( .INP(n81), .ZN(n79) );
  INVX0 U85 ( .INP(n77), .ZN(n75) );
  INVX0 U86 ( .INP(n81), .ZN(n80) );
  INVX0 U87 ( .INP(n81), .ZN(n78) );
  NBUFFX2 U88 ( .INP(n112), .Z(n57) );
  NBUFFX2 U89 ( .INP(n113), .Z(n61) );
  NBUFFX2 U90 ( .INP(n113), .Z(n60) );
  NBUFFX2 U91 ( .INP(n113), .Z(n59) );
  NBUFFX2 U92 ( .INP(n118), .Z(n63) );
  NBUFFX2 U93 ( .INP(n112), .Z(n58) );
  NBUFFX2 U94 ( .INP(n111), .Z(n54) );
  NBUFFX2 U95 ( .INP(n111), .Z(n53) );
  NBUFFX2 U96 ( .INP(n111), .Z(n55) );
  NBUFFX2 U97 ( .INP(n111), .Z(n56) );
  NBUFFX2 U98 ( .INP(reset), .Z(n52) );
  AND4X1 U99 ( .IN1(add_sum[1]), .IN2(n296), .IN3(n318), .IN4(n240), .Q(n134)
         );
  NAND3X0 U100 ( .IN1(n446), .IN2(n457), .IN3(add_sum[11]), .QN(n343) );
  NAND3X0 U101 ( .IN1(n464), .IN2(n475), .IN3(add_sum[14]), .QN(n242) );
  NAND3X0 U102 ( .IN1(n477), .IN2(n478), .IN3(add_sum[15]), .QN(n245) );
  INVX0 U103 ( .INP(N424), .ZN(n70) );
  NOR4X0 U104 ( .IN1(n321), .IN2(n355), .IN3(n490), .IN4(add_sum[22]), .QN(
        n142) );
  NAND3X0 U105 ( .IN1(n485), .IN2(n486), .IN3(add_sum[19]), .QN(n255) );
  NAND3X0 U106 ( .IN1(n480), .IN2(n484), .IN3(add_sum[18]), .QN(n249) );
  NBUFFX2 U107 ( .INP(add_new_exponent[5]), .Z(n84) );
  INVX0 U108 ( .INP(N580), .ZN(n74) );
  NBUFFX2 U109 ( .INP(add_new_exponent[5]), .Z(n82) );
  NBUFFX2 U110 ( .INP(add_new_exponent[6]), .Z(n86) );
  NBUFFX2 U111 ( .INP(add_new_exponent[5]), .Z(n83) );
  NBUFFX2 U112 ( .INP(add_new_exponent[7]), .Z(n87) );
  NBUFFX4 U113 ( .INP(add_new_exponent[6]), .Z(n85) );
  INVX0 U115 ( .INP(product_shift[26]), .ZN(n50) );
  INVX0 U116 ( .INP(n50), .ZN(n51) );
  INVX0 U117 ( .INP(n67), .ZN(n66) );
  INVX0 U118 ( .INP(N340), .ZN(n67) );
  INVX0 U119 ( .INP(n70), .ZN(n68) );
  INVX0 U120 ( .INP(n70), .ZN(n69) );
  INVX0 U121 ( .INP(n74), .ZN(n71) );
  INVX0 U122 ( .INP(n74), .ZN(n72) );
  INVX0 U123 ( .INP(n74), .ZN(n73) );
  INVX0 U124 ( .INP(N841), .ZN(n77) );
  INVX0 U125 ( .INP(add_new_exponent[4]), .ZN(n81) );
  XNOR2X1 U126 ( .IN1(n87), .IN2(\sub_419/carry[7] ), .Q(N723) );
  OR2X1 U127 ( .IN1(n86), .IN2(\sub_419/carry[6] ), .Q(\sub_419/carry[7] ) );
  XNOR2X1 U128 ( .IN1(\sub_419/carry[6] ), .IN2(n85), .Q(N722) );
  OR2X1 U129 ( .IN1(n83), .IN2(\sub_419/carry[5] ), .Q(\sub_419/carry[6] ) );
  XNOR2X1 U130 ( .IN1(\sub_419/carry[5] ), .IN2(n82), .Q(N721) );
  OR2X1 U131 ( .IN1(n80), .IN2(\sub_419/carry[4] ), .Q(\sub_419/carry[5] ) );
  AND2X1 U132 ( .IN1(n73), .IN2(N841), .Q(\sub_419/carry[4] ) );
  XOR2X1 U133 ( .IN1(n75), .IN2(n71), .Q(N719) );
  XNOR2X1 U134 ( .IN1(add_new_exponent[7]), .IN2(\sub_451/carry[7] ), .Q(N786)
         );
  OR2X1 U135 ( .IN1(n86), .IN2(\sub_451/carry[6] ), .Q(\sub_451/carry[7] ) );
  XNOR2X1 U136 ( .IN1(\sub_451/carry[6] ), .IN2(n85), .Q(N785) );
  OR2X1 U137 ( .IN1(n83), .IN2(\sub_451/carry[5] ), .Q(\sub_451/carry[6] ) );
  XNOR2X1 U138 ( .IN1(\sub_451/carry[5] ), .IN2(n82), .Q(N784) );
  OR2X1 U139 ( .IN1(n80), .IN2(\sub_451/carry[4] ), .Q(\sub_451/carry[5] ) );
  XNOR2X1 U140 ( .IN1(\sub_451/carry[4] ), .IN2(n79), .Q(N783) );
  AND2X1 U141 ( .IN1(\sub_451/carry[3] ), .IN2(n76), .Q(\sub_451/carry[4] ) );
  AND2X1 U142 ( .IN1(n69), .IN2(n73), .Q(\sub_451/carry[3] ) );
  XNOR2X1 U143 ( .IN1(add_new_exponent[7]), .IN2(\sub_435/carry[7] ), .Q(N755)
         );
  OR2X1 U144 ( .IN1(n86), .IN2(\sub_435/carry[6] ), .Q(\sub_435/carry[7] ) );
  XNOR2X1 U145 ( .IN1(\sub_435/carry[6] ), .IN2(n85), .Q(N754) );
  OR2X1 U146 ( .IN1(n83), .IN2(\sub_435/carry[5] ), .Q(\sub_435/carry[6] ) );
  XNOR2X1 U147 ( .IN1(\sub_435/carry[5] ), .IN2(n82), .Q(N753) );
  OR2X1 U148 ( .IN1(n79), .IN2(\sub_435/carry[4] ), .Q(\sub_435/carry[5] ) );
  XNOR2X1 U149 ( .IN1(\sub_435/carry[4] ), .IN2(n79), .Q(N752) );
  AND2X1 U150 ( .IN1(\sub_435/carry[3] ), .IN2(n76), .Q(\sub_435/carry[4] ) );
  XOR2X1 U151 ( .IN1(n75), .IN2(\sub_435/carry[3] ), .Q(N751) );
  AND2X1 U152 ( .IN1(\sub_435/carry[2] ), .IN2(n73), .Q(\sub_435/carry[3] ) );
  XOR2X1 U153 ( .IN1(n71), .IN2(\sub_435/carry[2] ), .Q(N750) );
  OR2X1 U154 ( .IN1(n69), .IN2(n66), .Q(\sub_435/carry[2] ) );
  XNOR2X1 U155 ( .IN1(n65), .IN2(n68), .Q(N749) );
  XNOR2X1 U156 ( .IN1(add_new_exponent[7]), .IN2(\sub_467/carry[7] ), .Q(N816)
         );
  OR2X1 U157 ( .IN1(n86), .IN2(\sub_467/carry[6] ), .Q(\sub_467/carry[7] ) );
  XNOR2X1 U158 ( .IN1(\sub_467/carry[6] ), .IN2(n85), .Q(N815) );
  OR2X1 U159 ( .IN1(n83), .IN2(\sub_467/carry[5] ), .Q(\sub_467/carry[6] ) );
  XNOR2X1 U160 ( .IN1(\sub_467/carry[5] ), .IN2(n82), .Q(N814) );
  OR2X1 U161 ( .IN1(n80), .IN2(\sub_467/carry[4] ), .Q(\sub_467/carry[5] ) );
  AND2X1 U162 ( .IN1(\sub_467/carry[3] ), .IN2(n76), .Q(\sub_467/carry[4] ) );
  XOR2X1 U163 ( .IN1(n75), .IN2(\sub_467/carry[3] ), .Q(N812) );
  AND2X1 U164 ( .IN1(\sub_467/carry[2] ), .IN2(n73), .Q(\sub_467/carry[3] ) );
  XOR2X1 U165 ( .IN1(n71), .IN2(\sub_467/carry[2] ), .Q(N811) );
  AND2X1 U166 ( .IN1(n66), .IN2(n69), .Q(\sub_467/carry[2] ) );
  XOR2X1 U167 ( .IN1(n68), .IN2(n65), .Q(N810) );
  XNOR2X1 U168 ( .IN1(add_new_exponent[7]), .IN2(\sub_499/carry[7] ), .Q(N873)
         );
  OR2X1 U169 ( .IN1(n86), .IN2(\sub_499/carry[6] ), .Q(\sub_499/carry[7] ) );
  XNOR2X1 U170 ( .IN1(\sub_499/carry[6] ), .IN2(n85), .Q(N872) );
  OR2X1 U171 ( .IN1(n83), .IN2(\sub_499/carry[5] ), .Q(\sub_499/carry[6] ) );
  XNOR2X1 U172 ( .IN1(\sub_499/carry[5] ), .IN2(n82), .Q(N871) );
  AND2X1 U173 ( .IN1(\sub_499/carry[4] ), .IN2(n80), .Q(\sub_499/carry[5] ) );
  XOR2X1 U174 ( .IN1(n78), .IN2(\sub_499/carry[4] ), .Q(N870) );
  OR2X1 U175 ( .IN1(N841), .IN2(\sub_499/carry[3] ), .Q(\sub_499/carry[4] ) );
  XNOR2X1 U176 ( .IN1(\sub_499/carry[3] ), .IN2(n76), .Q(N869) );
  OR2X1 U177 ( .IN1(n72), .IN2(\sub_499/carry[2] ), .Q(\sub_499/carry[3] ) );
  XNOR2X1 U178 ( .IN1(\sub_499/carry[2] ), .IN2(n72), .Q(N868) );
  OR2X1 U179 ( .IN1(n69), .IN2(n66), .Q(\sub_499/carry[2] ) );
  XNOR2X1 U180 ( .IN1(n65), .IN2(n68), .Q(N867) );
  XNOR2X1 U181 ( .IN1(n87), .IN2(\sub_483/carry[7] ), .Q(N845) );
  OR2X1 U182 ( .IN1(n86), .IN2(\sub_483/carry[6] ), .Q(\sub_483/carry[7] ) );
  XNOR2X1 U183 ( .IN1(\sub_483/carry[6] ), .IN2(n85), .Q(N844) );
  OR2X1 U184 ( .IN1(n83), .IN2(n79), .Q(\sub_483/carry[6] ) );
  XNOR2X1 U185 ( .IN1(n80), .IN2(n82), .Q(N843) );
  XNOR2X1 U186 ( .IN1(add_new_exponent[7]), .IN2(\sub_515/carry[7] ), .Q(N900)
         );
  OR2X1 U187 ( .IN1(n86), .IN2(\sub_515/carry[6] ), .Q(\sub_515/carry[7] ) );
  XNOR2X1 U188 ( .IN1(\sub_515/carry[6] ), .IN2(n85), .Q(N899) );
  OR2X1 U189 ( .IN1(n83), .IN2(\sub_515/carry[5] ), .Q(\sub_515/carry[6] ) );
  XNOR2X1 U190 ( .IN1(\sub_515/carry[5] ), .IN2(n82), .Q(N898) );
  AND2X1 U191 ( .IN1(\sub_515/carry[4] ), .IN2(n80), .Q(\sub_515/carry[5] ) );
  XOR2X1 U192 ( .IN1(n78), .IN2(\sub_515/carry[4] ), .Q(N897) );
  OR2X1 U193 ( .IN1(n75), .IN2(\sub_515/carry[3] ), .Q(\sub_515/carry[4] ) );
  XNOR2X1 U194 ( .IN1(\sub_515/carry[3] ), .IN2(n76), .Q(N896) );
  OR2X1 U195 ( .IN1(n72), .IN2(n69), .Q(\sub_515/carry[3] ) );
  XNOR2X1 U196 ( .IN1(n68), .IN2(n72), .Q(N895) );
  XNOR2X1 U197 ( .IN1(add_new_exponent[7]), .IN2(\sub_547/carry[7] ), .Q(N951)
         );
  OR2X1 U198 ( .IN1(n86), .IN2(\sub_547/carry[6] ), .Q(\sub_547/carry[7] ) );
  XNOR2X1 U199 ( .IN1(\sub_547/carry[6] ), .IN2(n85), .Q(N950) );
  OR2X1 U200 ( .IN1(n83), .IN2(\sub_547/carry[5] ), .Q(\sub_547/carry[6] ) );
  XNOR2X1 U201 ( .IN1(\sub_547/carry[5] ), .IN2(n84), .Q(N949) );
  AND2X1 U202 ( .IN1(\sub_547/carry[4] ), .IN2(n78), .Q(\sub_547/carry[5] ) );
  OR2X1 U203 ( .IN1(n76), .IN2(n72), .Q(\sub_547/carry[4] ) );
  XNOR2X1 U204 ( .IN1(n73), .IN2(n76), .Q(N947) );
  XNOR2X1 U205 ( .IN1(add_new_exponent[7]), .IN2(\sub_531/carry[7] ), .Q(N926)
         );
  OR2X1 U206 ( .IN1(n85), .IN2(\sub_531/carry[6] ), .Q(\sub_531/carry[7] ) );
  XNOR2X1 U207 ( .IN1(\sub_531/carry[6] ), .IN2(n85), .Q(N925) );
  OR2X1 U208 ( .IN1(n82), .IN2(\sub_531/carry[5] ), .Q(\sub_531/carry[6] ) );
  XNOR2X1 U209 ( .IN1(\sub_531/carry[5] ), .IN2(n84), .Q(N924) );
  AND2X1 U210 ( .IN1(\sub_531/carry[4] ), .IN2(n80), .Q(\sub_531/carry[5] ) );
  OR2X1 U211 ( .IN1(n76), .IN2(\sub_531/carry[3] ), .Q(\sub_531/carry[4] ) );
  XNOR2X1 U212 ( .IN1(\sub_531/carry[3] ), .IN2(n76), .Q(N922) );
  OR2X1 U213 ( .IN1(n72), .IN2(\sub_531/carry[2] ), .Q(\sub_531/carry[3] ) );
  XNOR2X1 U214 ( .IN1(\sub_531/carry[2] ), .IN2(n72), .Q(N921) );
  AND2X1 U215 ( .IN1(n66), .IN2(n69), .Q(\sub_531/carry[2] ) );
  XOR2X1 U216 ( .IN1(n68), .IN2(n66), .Q(N920) );
  XNOR2X1 U217 ( .IN1(add_new_exponent[7]), .IN2(\sub_563/carry[7] ), .Q(N975)
         );
  OR2X1 U218 ( .IN1(n85), .IN2(\sub_563/carry[6] ), .Q(\sub_563/carry[7] ) );
  XNOR2X1 U219 ( .IN1(\sub_563/carry[6] ), .IN2(n85), .Q(N974) );
  OR2X1 U220 ( .IN1(n82), .IN2(\sub_563/carry[5] ), .Q(\sub_563/carry[6] ) );
  XNOR2X1 U221 ( .IN1(\sub_563/carry[5] ), .IN2(add_new_exponent[5]), .Q(N973)
         );
  AND2X1 U222 ( .IN1(\sub_563/carry[4] ), .IN2(n80), .Q(\sub_563/carry[5] ) );
  XOR2X1 U223 ( .IN1(n78), .IN2(\sub_563/carry[4] ), .Q(N972) );
  OR2X1 U224 ( .IN1(n76), .IN2(\sub_563/carry[3] ), .Q(\sub_563/carry[4] ) );
  XNOR2X1 U225 ( .IN1(\sub_563/carry[3] ), .IN2(n76), .Q(N971) );
  AND2X1 U226 ( .IN1(\sub_563/carry[2] ), .IN2(n73), .Q(\sub_563/carry[3] ) );
  XOR2X1 U227 ( .IN1(n71), .IN2(\sub_563/carry[2] ), .Q(N970) );
  OR2X1 U228 ( .IN1(n68), .IN2(N340), .Q(\sub_563/carry[2] ) );
  XNOR2X1 U229 ( .IN1(n65), .IN2(n69), .Q(N969) );
  XNOR2X1 U230 ( .IN1(n87), .IN2(\sub_595/carry[7] ), .Q(N1020) );
  OR2X1 U231 ( .IN1(n85), .IN2(\sub_595/carry[6] ), .Q(\sub_595/carry[7] ) );
  XNOR2X1 U232 ( .IN1(\sub_595/carry[6] ), .IN2(n85), .Q(N1019) );
  OR2X1 U233 ( .IN1(n82), .IN2(\sub_595/carry[5] ), .Q(\sub_595/carry[6] ) );
  XNOR2X1 U234 ( .IN1(\sub_595/carry[5] ), .IN2(n84), .Q(N1018) );
  AND2X1 U235 ( .IN1(\sub_595/carry[4] ), .IN2(n80), .Q(\sub_595/carry[5] ) );
  XOR2X1 U236 ( .IN1(n78), .IN2(\sub_595/carry[4] ), .Q(N1017) );
  OR2X1 U237 ( .IN1(n76), .IN2(\sub_595/carry[3] ), .Q(\sub_595/carry[4] ) );
  XNOR2X1 U238 ( .IN1(\sub_595/carry[3] ), .IN2(n76), .Q(N1016) );
  AND2X1 U239 ( .IN1(\sub_595/carry[2] ), .IN2(n73), .Q(\sub_595/carry[3] ) );
  XOR2X1 U240 ( .IN1(n71), .IN2(\sub_595/carry[2] ), .Q(N1015) );
  AND2X1 U241 ( .IN1(n66), .IN2(n69), .Q(\sub_595/carry[2] ) );
  XOR2X1 U242 ( .IN1(n68), .IN2(n66), .Q(N1014) );
  XNOR2X1 U243 ( .IN1(n87), .IN2(\sub_579/carry[7] ), .Q(N998) );
  OR2X1 U244 ( .IN1(n85), .IN2(\sub_579/carry[6] ), .Q(\sub_579/carry[7] ) );
  XNOR2X1 U245 ( .IN1(\sub_579/carry[6] ), .IN2(n85), .Q(N997) );
  OR2X1 U246 ( .IN1(n82), .IN2(\sub_579/carry[5] ), .Q(\sub_579/carry[6] ) );
  XNOR2X1 U247 ( .IN1(\sub_579/carry[5] ), .IN2(n84), .Q(N996) );
  AND2X1 U248 ( .IN1(\sub_579/carry[4] ), .IN2(n80), .Q(\sub_579/carry[5] ) );
  XOR2X1 U249 ( .IN1(n78), .IN2(\sub_579/carry[4] ), .Q(N995) );
  OR2X1 U250 ( .IN1(n76), .IN2(\sub_579/carry[3] ), .Q(\sub_579/carry[4] ) );
  XNOR2X1 U251 ( .IN1(\sub_579/carry[3] ), .IN2(n76), .Q(N994) );
  AND2X1 U252 ( .IN1(n69), .IN2(n73), .Q(\sub_579/carry[3] ) );
  XNOR2X1 U253 ( .IN1(n87), .IN2(\sub_259/carry[7] ), .Q(N347) );
  OR2X1 U254 ( .IN1(n85), .IN2(\sub_259/carry[6] ), .Q(\sub_259/carry[7] ) );
  XNOR2X1 U255 ( .IN1(\sub_259/carry[6] ), .IN2(n85), .Q(N346) );
  OR2X1 U256 ( .IN1(n82), .IN2(\sub_259/carry[5] ), .Q(\sub_259/carry[6] ) );
  XNOR2X1 U257 ( .IN1(\sub_259/carry[5] ), .IN2(n84), .Q(N345) );
  OR2X1 U258 ( .IN1(n79), .IN2(\sub_259/carry[4] ), .Q(\sub_259/carry[5] ) );
  XNOR2X1 U259 ( .IN1(\sub_259/carry[4] ), .IN2(n79), .Q(N344) );
  OR2X1 U260 ( .IN1(n76), .IN2(\sub_259/carry[3] ), .Q(\sub_259/carry[4] ) );
  XNOR2X1 U261 ( .IN1(\sub_259/carry[3] ), .IN2(n76), .Q(N343) );
  OR2X1 U262 ( .IN1(n72), .IN2(N424), .Q(\sub_259/carry[3] ) );
  XNOR2X1 U263 ( .IN1(n68), .IN2(n72), .Q(N342) );
  XNOR2X1 U264 ( .IN1(n87), .IN2(\sub_291/carry[7] ), .Q(N430) );
  OR2X1 U265 ( .IN1(n85), .IN2(\sub_291/carry[6] ), .Q(\sub_291/carry[7] ) );
  XNOR2X1 U266 ( .IN1(\sub_291/carry[6] ), .IN2(n85), .Q(N429) );
  OR2X1 U267 ( .IN1(n82), .IN2(\sub_291/carry[5] ), .Q(\sub_291/carry[6] ) );
  XNOR2X1 U268 ( .IN1(\sub_291/carry[5] ), .IN2(n84), .Q(N428) );
  OR2X1 U269 ( .IN1(n79), .IN2(\sub_291/carry[4] ), .Q(\sub_291/carry[5] ) );
  XNOR2X1 U270 ( .IN1(\sub_291/carry[4] ), .IN2(n78), .Q(N427) );
  OR2X1 U271 ( .IN1(n76), .IN2(n72), .Q(\sub_291/carry[4] ) );
  XNOR2X1 U272 ( .IN1(n87), .IN2(\sub_307/carry[7] ), .Q(N470) );
  OR2X1 U273 ( .IN1(n85), .IN2(\sub_307/carry[6] ), .Q(\sub_307/carry[7] ) );
  XNOR2X1 U274 ( .IN1(\sub_307/carry[6] ), .IN2(n85), .Q(N469) );
  OR2X1 U275 ( .IN1(n82), .IN2(\sub_307/carry[5] ), .Q(\sub_307/carry[6] ) );
  XNOR2X1 U276 ( .IN1(\sub_307/carry[5] ), .IN2(n84), .Q(N468) );
  OR2X1 U277 ( .IN1(n79), .IN2(\sub_307/carry[4] ), .Q(\sub_307/carry[5] ) );
  XNOR2X1 U278 ( .IN1(\sub_307/carry[4] ), .IN2(n79), .Q(N467) );
  OR2X1 U279 ( .IN1(n76), .IN2(\sub_307/carry[3] ), .Q(\sub_307/carry[4] ) );
  XNOR2X1 U280 ( .IN1(\sub_307/carry[3] ), .IN2(n75), .Q(N466) );
  AND2X1 U281 ( .IN1(\sub_307/carry[2] ), .IN2(n73), .Q(\sub_307/carry[3] ) );
  XOR2X1 U282 ( .IN1(n71), .IN2(\sub_307/carry[2] ), .Q(N465) );
  OR2X1 U283 ( .IN1(N424), .IN2(N340), .Q(\sub_307/carry[2] ) );
  XNOR2X1 U284 ( .IN1(n65), .IN2(n69), .Q(N464) );
  XNOR2X1 U285 ( .IN1(n87), .IN2(\sub_275/carry[7] ), .Q(N389) );
  OR2X1 U286 ( .IN1(n86), .IN2(\sub_275/carry[6] ), .Q(\sub_275/carry[7] ) );
  XNOR2X1 U287 ( .IN1(\sub_275/carry[6] ), .IN2(n85), .Q(N388) );
  OR2X1 U288 ( .IN1(n83), .IN2(\sub_275/carry[5] ), .Q(\sub_275/carry[6] ) );
  XNOR2X1 U289 ( .IN1(\sub_275/carry[5] ), .IN2(n84), .Q(N387) );
  OR2X1 U290 ( .IN1(n79), .IN2(\sub_275/carry[4] ), .Q(\sub_275/carry[5] ) );
  XNOR2X1 U291 ( .IN1(\sub_275/carry[4] ), .IN2(n78), .Q(N386) );
  OR2X1 U292 ( .IN1(n76), .IN2(\sub_275/carry[3] ), .Q(\sub_275/carry[4] ) );
  XNOR2X1 U293 ( .IN1(\sub_275/carry[3] ), .IN2(n75), .Q(N385) );
  OR2X1 U294 ( .IN1(n72), .IN2(\sub_275/carry[2] ), .Q(\sub_275/carry[3] ) );
  XNOR2X1 U295 ( .IN1(\sub_275/carry[2] ), .IN2(n72), .Q(N384) );
  AND2X1 U296 ( .IN1(n66), .IN2(n69), .Q(\sub_275/carry[2] ) );
  XOR2X1 U297 ( .IN1(n68), .IN2(n65), .Q(N383) );
  XNOR2X1 U298 ( .IN1(n87), .IN2(\sub_323/carry[7] ), .Q(N509) );
  OR2X1 U299 ( .IN1(n86), .IN2(\sub_323/carry[6] ), .Q(\sub_323/carry[7] ) );
  XNOR2X1 U300 ( .IN1(\sub_323/carry[6] ), .IN2(n85), .Q(N508) );
  OR2X1 U301 ( .IN1(n83), .IN2(\sub_323/carry[5] ), .Q(\sub_323/carry[6] ) );
  XNOR2X1 U302 ( .IN1(\sub_323/carry[5] ), .IN2(n84), .Q(N507) );
  OR2X1 U303 ( .IN1(n80), .IN2(\sub_323/carry[4] ), .Q(\sub_323/carry[5] ) );
  XNOR2X1 U304 ( .IN1(\sub_323/carry[4] ), .IN2(n78), .Q(N506) );
  OR2X1 U305 ( .IN1(n75), .IN2(\sub_323/carry[3] ), .Q(\sub_323/carry[4] ) );
  XNOR2X1 U306 ( .IN1(\sub_323/carry[3] ), .IN2(n75), .Q(N505) );
  AND2X1 U307 ( .IN1(n69), .IN2(n73), .Q(\sub_323/carry[3] ) );
  XOR2X1 U308 ( .IN1(n71), .IN2(n68), .Q(N504) );
  XNOR2X1 U309 ( .IN1(n87), .IN2(\sub_355/carry[7] ), .Q(N585) );
  OR2X1 U310 ( .IN1(n86), .IN2(\sub_355/carry[6] ), .Q(\sub_355/carry[7] ) );
  XNOR2X1 U311 ( .IN1(\sub_355/carry[6] ), .IN2(n85), .Q(N584) );
  OR2X1 U312 ( .IN1(n83), .IN2(\sub_355/carry[5] ), .Q(\sub_355/carry[6] ) );
  XNOR2X1 U313 ( .IN1(\sub_355/carry[5] ), .IN2(n84), .Q(N583) );
  OR2X1 U314 ( .IN1(n79), .IN2(n76), .Q(\sub_355/carry[5] ) );
  XNOR2X1 U315 ( .IN1(N841), .IN2(n79), .Q(N582) );
  XNOR2X1 U316 ( .IN1(n87), .IN2(\sub_339/carry[7] ), .Q(N547) );
  OR2X1 U317 ( .IN1(n86), .IN2(\sub_339/carry[6] ), .Q(\sub_339/carry[7] ) );
  XNOR2X1 U318 ( .IN1(\sub_339/carry[6] ), .IN2(n85), .Q(N546) );
  OR2X1 U319 ( .IN1(n83), .IN2(\sub_339/carry[5] ), .Q(\sub_339/carry[6] ) );
  XNOR2X1 U320 ( .IN1(\sub_339/carry[5] ), .IN2(n82), .Q(N545) );
  OR2X1 U321 ( .IN1(n80), .IN2(\sub_339/carry[4] ), .Q(\sub_339/carry[5] ) );
  XNOR2X1 U322 ( .IN1(\sub_339/carry[4] ), .IN2(n79), .Q(N544) );
  OR2X1 U323 ( .IN1(n76), .IN2(\sub_339/carry[3] ), .Q(\sub_339/carry[4] ) );
  XNOR2X1 U324 ( .IN1(\sub_339/carry[3] ), .IN2(n75), .Q(N543) );
  AND2X1 U325 ( .IN1(\sub_339/carry[2] ), .IN2(n73), .Q(\sub_339/carry[3] ) );
  XOR2X1 U326 ( .IN1(n71), .IN2(\sub_339/carry[2] ), .Q(N542) );
  AND2X1 U327 ( .IN1(n66), .IN2(n69), .Q(\sub_339/carry[2] ) );
  XOR2X1 U328 ( .IN1(n68), .IN2(N340), .Q(N541) );
  XNOR2X1 U329 ( .IN1(n87), .IN2(\sub_387/carry[7] ), .Q(N656) );
  OR2X1 U330 ( .IN1(n86), .IN2(\sub_387/carry[6] ), .Q(\sub_387/carry[7] ) );
  XNOR2X1 U331 ( .IN1(\sub_387/carry[6] ), .IN2(n85), .Q(N655) );
  OR2X1 U332 ( .IN1(n83), .IN2(\sub_387/carry[5] ), .Q(\sub_387/carry[6] ) );
  XNOR2X1 U333 ( .IN1(\sub_387/carry[5] ), .IN2(n84), .Q(N654) );
  OR2X1 U334 ( .IN1(n80), .IN2(\sub_387/carry[4] ), .Q(\sub_387/carry[5] ) );
  XNOR2X1 U335 ( .IN1(\sub_387/carry[4] ), .IN2(n78), .Q(N653) );
  AND2X1 U336 ( .IN1(\sub_387/carry[3] ), .IN2(n76), .Q(\sub_387/carry[4] ) );
  OR2X1 U337 ( .IN1(n72), .IN2(n68), .Q(\sub_387/carry[3] ) );
  XNOR2X1 U338 ( .IN1(N424), .IN2(n72), .Q(N651) );
  XNOR2X1 U339 ( .IN1(n87), .IN2(\sub_403/carry[7] ), .Q(N690) );
  OR2X1 U340 ( .IN1(n86), .IN2(\sub_403/carry[6] ), .Q(\sub_403/carry[7] ) );
  XNOR2X1 U341 ( .IN1(\sub_403/carry[6] ), .IN2(n85), .Q(N689) );
  OR2X1 U342 ( .IN1(n83), .IN2(\sub_403/carry[5] ), .Q(\sub_403/carry[6] ) );
  XNOR2X1 U343 ( .IN1(\sub_403/carry[5] ), .IN2(n84), .Q(N688) );
  OR2X1 U344 ( .IN1(n80), .IN2(\sub_403/carry[4] ), .Q(\sub_403/carry[5] ) );
  XNOR2X1 U345 ( .IN1(\sub_403/carry[4] ), .IN2(n79), .Q(N687) );
  AND2X1 U346 ( .IN1(\sub_403/carry[3] ), .IN2(n76), .Q(\sub_403/carry[4] ) );
  XOR2X1 U347 ( .IN1(n75), .IN2(\sub_403/carry[3] ), .Q(N686) );
  OR2X1 U348 ( .IN1(n72), .IN2(\sub_403/carry[2] ), .Q(\sub_403/carry[3] ) );
  XNOR2X1 U349 ( .IN1(\sub_403/carry[2] ), .IN2(n71), .Q(N685) );
  AND2X1 U350 ( .IN1(n66), .IN2(n69), .Q(\sub_403/carry[2] ) );
  XOR2X1 U351 ( .IN1(n68), .IN2(N340), .Q(N684) );
  XNOR2X1 U352 ( .IN1(n87), .IN2(\sub_371/carry[7] ), .Q(N621) );
  OR2X1 U353 ( .IN1(n86), .IN2(\sub_371/carry[6] ), .Q(\sub_371/carry[7] ) );
  XNOR2X1 U354 ( .IN1(\sub_371/carry[6] ), .IN2(n85), .Q(N620) );
  OR2X1 U355 ( .IN1(n83), .IN2(\sub_371/carry[5] ), .Q(\sub_371/carry[6] ) );
  XNOR2X1 U356 ( .IN1(\sub_371/carry[5] ), .IN2(n84), .Q(N619) );
  OR2X1 U357 ( .IN1(n80), .IN2(\sub_371/carry[4] ), .Q(\sub_371/carry[5] ) );
  XNOR2X1 U358 ( .IN1(\sub_371/carry[4] ), .IN2(n78), .Q(N618) );
  AND2X1 U359 ( .IN1(\sub_371/carry[3] ), .IN2(n76), .Q(\sub_371/carry[4] ) );
  XOR2X1 U360 ( .IN1(n75), .IN2(\sub_371/carry[3] ), .Q(N617) );
  OR2X1 U361 ( .IN1(n72), .IN2(\sub_371/carry[2] ), .Q(\sub_371/carry[3] ) );
  XNOR2X1 U362 ( .IN1(\sub_371/carry[2] ), .IN2(n71), .Q(N616) );
  XNOR2X1 U363 ( .IN1(n65), .IN2(n68), .Q(N615) );
  NOR2X0 U364 ( .IN1(n69), .IN2(n65), .QN(n101) );
  AO21X1 U365 ( .IN1(n69), .IN2(n66), .IN3(n101), .Q(N298) );
  NOR2X0 U366 ( .IN1(\sub_307/carry[2] ), .IN2(n73), .QN(n102) );
  AO21X1 U367 ( .IN1(n73), .IN2(\sub_563/carry[2] ), .IN3(n102), .Q(N299) );
  NOR2X0 U368 ( .IN1(n107), .IN2(n75), .QN(n103) );
  AO21X1 U369 ( .IN1(n76), .IN2(n107), .IN3(n103), .Q(N300) );
  NOR2X0 U370 ( .IN1(n108), .IN2(n80), .QN(n104) );
  AO21X1 U371 ( .IN1(n80), .IN2(n108), .IN3(n104), .Q(N301) );
  NOR2X0 U372 ( .IN1(n109), .IN2(n83), .QN(n105) );
  AO21X1 U373 ( .IN1(n84), .IN2(n109), .IN3(n105), .Q(N302) );
  XNOR2X1 U374 ( .IN1(n86), .IN2(n110), .Q(N303) );
  NOR2X0 U375 ( .IN1(n86), .IN2(n110), .QN(n106) );
  XOR2X1 U376 ( .IN1(n87), .IN2(n106), .Q(N304) );
  AO222X1 U377 ( .IN1(N133), .IN2(n53), .IN3(product_shift[9]), .IN4(n57), 
        .IN5(N82), .IN6(n59), .Q(product2[9]) );
  AO222X1 U378 ( .IN1(N132), .IN2(n53), .IN3(product_shift[8]), .IN4(n58), 
        .IN5(N81), .IN6(n59), .Q(product2[8]) );
  AO222X1 U379 ( .IN1(N131), .IN2(n53), .IN3(product_shift[7]), .IN4(n58), 
        .IN5(N80), .IN6(n59), .Q(product2[7]) );
  AO222X1 U380 ( .IN1(N130), .IN2(n53), .IN3(product_shift[6]), .IN4(n58), 
        .IN5(N79), .IN6(n59), .Q(product2[6]) );
  AO222X1 U381 ( .IN1(N129), .IN2(n53), .IN3(product_shift[5]), .IN4(n58), 
        .IN5(N78), .IN6(n59), .Q(product2[5]) );
  AO222X1 U382 ( .IN1(N174), .IN2(n53), .IN3(product_shift[49]), .IN4(n58), 
        .IN5(n59), .IN6(N123), .Q(product2[50]) );
  AO222X1 U383 ( .IN1(N128), .IN2(n53), .IN3(product_shift[4]), .IN4(n58), 
        .IN5(N77), .IN6(n59), .Q(product2[4]) );
  AO222X1 U384 ( .IN1(N173), .IN2(n53), .IN3(product_shift[49]), .IN4(n58), 
        .IN5(N122), .IN6(n59), .Q(product2[49]) );
  AO222X1 U385 ( .IN1(N172), .IN2(n53), .IN3(product_shift[48]), .IN4(n58), 
        .IN5(N121), .IN6(n59), .Q(product2[48]) );
  AO222X1 U386 ( .IN1(N171), .IN2(n53), .IN3(product_shift[47]), .IN4(n58), 
        .IN5(N120), .IN6(n59), .Q(product2[47]) );
  AO222X1 U387 ( .IN1(N170), .IN2(n53), .IN3(product_shift[46]), .IN4(n58), 
        .IN5(N119), .IN6(n59), .Q(product2[46]) );
  AO222X1 U388 ( .IN1(N169), .IN2(n53), .IN3(product_shift[45]), .IN4(n58), 
        .IN5(N118), .IN6(n59), .Q(product2[45]) );
  AO222X1 U389 ( .IN1(N168), .IN2(n54), .IN3(product_shift[44]), .IN4(n58), 
        .IN5(N117), .IN6(n60), .Q(product2[44]) );
  AO222X1 U390 ( .IN1(N167), .IN2(n54), .IN3(product_shift[43]), .IN4(n57), 
        .IN5(N116), .IN6(n60), .Q(product2[43]) );
  AO222X1 U391 ( .IN1(N166), .IN2(n54), .IN3(product_shift[42]), .IN4(n58), 
        .IN5(N115), .IN6(n60), .Q(product2[42]) );
  AO222X1 U392 ( .IN1(N165), .IN2(n54), .IN3(product_shift[41]), .IN4(n112), 
        .IN5(N114), .IN6(n60), .Q(product2[41]) );
  AO222X1 U393 ( .IN1(N164), .IN2(n54), .IN3(product_shift[40]), .IN4(n112), 
        .IN5(N113), .IN6(n60), .Q(product2[40]) );
  AO222X1 U394 ( .IN1(N127), .IN2(n54), .IN3(product_shift[3]), .IN4(n112), 
        .IN5(N76), .IN6(n60), .Q(product2[3]) );
  AO222X1 U395 ( .IN1(N163), .IN2(n54), .IN3(product_shift[39]), .IN4(n112), 
        .IN5(N112), .IN6(n60), .Q(product2[39]) );
  AO222X1 U396 ( .IN1(N162), .IN2(n54), .IN3(product_shift[38]), .IN4(n112), 
        .IN5(N111), .IN6(n60), .Q(product2[38]) );
  AO222X1 U397 ( .IN1(N161), .IN2(n54), .IN3(product_shift[37]), .IN4(n112), 
        .IN5(N110), .IN6(n60), .Q(product2[37]) );
  AO222X1 U398 ( .IN1(N160), .IN2(n54), .IN3(product_shift[36]), .IN4(n112), 
        .IN5(N109), .IN6(n60), .Q(product2[36]) );
  AO222X1 U399 ( .IN1(N159), .IN2(n54), .IN3(product_shift[35]), .IN4(n112), 
        .IN5(N108), .IN6(n60), .Q(product2[35]) );
  AO222X1 U400 ( .IN1(N158), .IN2(n54), .IN3(n6), .IN4(n112), .IN5(N107), 
        .IN6(n60), .Q(product2[34]) );
  AO222X1 U401 ( .IN1(N157), .IN2(n55), .IN3(n12), .IN4(n112), .IN5(N106), 
        .IN6(n113), .Q(product2[33]) );
  AO222X1 U402 ( .IN1(N156), .IN2(n55), .IN3(n18), .IN4(n58), .IN5(N105), 
        .IN6(n113), .Q(product2[32]) );
  AO222X1 U403 ( .IN1(N155), .IN2(n55), .IN3(n24), .IN4(n112), .IN5(N104), 
        .IN6(n113), .Q(product2[31]) );
  AO222X1 U404 ( .IN1(N154), .IN2(n55), .IN3(n30), .IN4(n57), .IN5(N103), 
        .IN6(n113), .Q(product2[30]) );
  AO222X1 U405 ( .IN1(N126), .IN2(n55), .IN3(product_shift[2]), .IN4(n112), 
        .IN5(N75), .IN6(n113), .Q(product2[2]) );
  AO222X1 U406 ( .IN1(N153), .IN2(n55), .IN3(n36), .IN4(n112), .IN5(N102), 
        .IN6(n113), .Q(product2[29]) );
  AO222X1 U407 ( .IN1(N152), .IN2(n55), .IN3(n42), .IN4(n112), .IN5(N101), 
        .IN6(n113), .Q(product2[28]) );
  AO222X1 U408 ( .IN1(N151), .IN2(n55), .IN3(n49), .IN4(n112), .IN5(N100), 
        .IN6(n113), .Q(product2[27]) );
  AO222X1 U409 ( .IN1(N150), .IN2(n55), .IN3(n51), .IN4(n112), .IN5(N99), 
        .IN6(n113), .Q(product2[26]) );
  AO222X1 U410 ( .IN1(N149), .IN2(n55), .IN3(product_shift[25]), .IN4(n112), 
        .IN5(N98), .IN6(n113), .Q(product2[25]) );
  AO222X1 U411 ( .IN1(N148), .IN2(n55), .IN3(product_shift[24]), .IN4(n112), 
        .IN5(N97), .IN6(n59), .Q(product2[24]) );
  AO222X1 U412 ( .IN1(N146), .IN2(n54), .IN3(product_shift[22]), .IN4(n58), 
        .IN5(N95), .IN6(n61), .Q(product2[22]) );
  AO222X1 U413 ( .IN1(N145), .IN2(n56), .IN3(product_shift[21]), .IN4(n57), 
        .IN5(N94), .IN6(n61), .Q(product2[21]) );
  AO222X1 U414 ( .IN1(N144), .IN2(n55), .IN3(product_shift[20]), .IN4(n57), 
        .IN5(N93), .IN6(n61), .Q(product2[20]) );
  AO222X1 U415 ( .IN1(N125), .IN2(n56), .IN3(n57), .IN4(product_shift[1]), 
        .IN5(N74), .IN6(n61), .Q(product2[1]) );
  AO222X1 U416 ( .IN1(N143), .IN2(n56), .IN3(product_shift[19]), .IN4(n57), 
        .IN5(N92), .IN6(n61), .Q(product2[19]) );
  AO222X1 U417 ( .IN1(N142), .IN2(n56), .IN3(product_shift[18]), .IN4(n57), 
        .IN5(N91), .IN6(n61), .Q(product2[18]) );
  AO222X1 U418 ( .IN1(N141), .IN2(n56), .IN3(product_shift[17]), .IN4(n57), 
        .IN5(N90), .IN6(n61), .Q(product2[17]) );
  AO222X1 U419 ( .IN1(N140), .IN2(n56), .IN3(product_shift[16]), .IN4(n57), 
        .IN5(N89), .IN6(n61), .Q(product2[16]) );
  AO222X1 U420 ( .IN1(N139), .IN2(n56), .IN3(product_shift[15]), .IN4(n57), 
        .IN5(N88), .IN6(n61), .Q(product2[15]) );
  AO222X1 U421 ( .IN1(N138), .IN2(n56), .IN3(product_shift[14]), .IN4(n57), 
        .IN5(N87), .IN6(n61), .Q(product2[14]) );
  AO222X1 U422 ( .IN1(N137), .IN2(n56), .IN3(product_shift[13]), .IN4(n57), 
        .IN5(N86), .IN6(n61), .Q(product2[13]) );
  AO222X1 U423 ( .IN1(N136), .IN2(n56), .IN3(product_shift[12]), .IN4(n57), 
        .IN5(N85), .IN6(n61), .Q(product2[12]) );
  AO222X1 U424 ( .IN1(N135), .IN2(n56), .IN3(product_shift[11]), .IN4(n57), 
        .IN5(N84), .IN6(n60), .Q(product2[11]) );
  AO222X1 U425 ( .IN1(N134), .IN2(n56), .IN3(product_shift[10]), .IN4(n58), 
        .IN5(N83), .IN6(n61), .Q(product2[10]) );
  AND2X1 U426 ( .IN1(product_shift[0]), .IN2(n114), .Q(n113) );
  XNOR2X1 U427 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n112) );
  NOR2X0 U428 ( .IN1(n114), .IN2(product_shift[0]), .QN(n111) );
  INVX0 U429 ( .INP(product_shift[1]), .ZN(n114) );
  AO222X1 U430 ( .IN1(N199), .IN2(n115), .IN3(n62), .IN4(n117), .IN5(n118), 
        .IN6(add_new_exponent[7]), .Q(add_updated_exponent[7]) );
  NAND2X0 U431 ( .IN1(n119), .IN2(n120), .QN(n117) );
  NOR4X0 U432 ( .IN1(n121), .IN2(n122), .IN3(n123), .IN4(n124), .QN(n120) );
  AO222X1 U433 ( .IN1(N755), .IN2(n125), .IN3(N786), .IN4(n126), .IN5(N723), 
        .IN6(n127), .Q(n124) );
  AO222X1 U434 ( .IN1(N845), .IN2(n128), .IN3(N873), .IN4(n129), .IN5(N816), 
        .IN6(n130), .Q(n123) );
  AO222X1 U435 ( .IN1(N926), .IN2(n131), .IN3(N951), .IN4(n132), .IN5(N900), 
        .IN6(n133), .Q(n122) );
  AO222X1 U436 ( .IN1(N998), .IN2(n134), .IN3(N1020), .IN4(n135), .IN5(N975), 
        .IN6(n136), .Q(n121) );
  NOR4X0 U437 ( .IN1(n137), .IN2(n138), .IN3(n139), .IN4(n140), .QN(n119) );
  AO222X1 U438 ( .IN1(N304), .IN2(n141), .IN3(N347), .IN4(n142), .IN5(
        add_sum[23]), .IN6(add_new_exponent[7]), .Q(n140) );
  AO222X1 U439 ( .IN1(N389), .IN2(n143), .IN3(N470), .IN4(n144), .IN5(N430), 
        .IN6(n145), .Q(n139) );
  AO222X1 U440 ( .IN1(N547), .IN2(n146), .IN3(N585), .IN4(n147), .IN5(N509), 
        .IN6(n148), .Q(n138) );
  AO222X1 U441 ( .IN1(N621), .IN2(n149), .IN3(N690), .IN4(n150), .IN5(N656), 
        .IN6(n151), .Q(n137) );
  AO222X1 U442 ( .IN1(N198), .IN2(n115), .IN3(n62), .IN4(n152), .IN5(
        add_new_exponent[6]), .IN6(n118), .Q(add_updated_exponent[6]) );
  NAND2X0 U443 ( .IN1(n153), .IN2(n154), .QN(n152) );
  NOR4X0 U444 ( .IN1(n155), .IN2(n156), .IN3(n157), .IN4(n158), .QN(n154) );
  AO222X1 U445 ( .IN1(N754), .IN2(n125), .IN3(N785), .IN4(n126), .IN5(N722), 
        .IN6(n127), .Q(n158) );
  AO222X1 U446 ( .IN1(N844), .IN2(n128), .IN3(N872), .IN4(n129), .IN5(N815), 
        .IN6(n130), .Q(n157) );
  AO222X1 U447 ( .IN1(N925), .IN2(n131), .IN3(N950), .IN4(n132), .IN5(N899), 
        .IN6(n133), .Q(n156) );
  AO222X1 U448 ( .IN1(N997), .IN2(n134), .IN3(N1019), .IN4(n135), .IN5(N974), 
        .IN6(n136), .Q(n155) );
  NOR4X0 U449 ( .IN1(n159), .IN2(n160), .IN3(n161), .IN4(n162), .QN(n153) );
  AO222X1 U450 ( .IN1(N303), .IN2(n141), .IN3(N346), .IN4(n142), .IN5(
        add_new_exponent[6]), .IN6(add_sum[23]), .Q(n162) );
  AO222X1 U451 ( .IN1(N388), .IN2(n143), .IN3(N469), .IN4(n144), .IN5(N429), 
        .IN6(n145), .Q(n161) );
  AO222X1 U452 ( .IN1(N546), .IN2(n146), .IN3(N584), .IN4(n147), .IN5(N508), 
        .IN6(n148), .Q(n160) );
  AO222X1 U453 ( .IN1(N620), .IN2(n149), .IN3(N689), .IN4(n150), .IN5(N655), 
        .IN6(n151), .Q(n159) );
  AO222X1 U454 ( .IN1(N197), .IN2(n115), .IN3(n62), .IN4(n163), .IN5(n83), 
        .IN6(n118), .Q(add_updated_exponent[5]) );
  NAND2X0 U455 ( .IN1(n164), .IN2(n165), .QN(n163) );
  NOR4X0 U456 ( .IN1(n166), .IN2(n167), .IN3(n168), .IN4(n169), .QN(n165) );
  AO222X1 U457 ( .IN1(N753), .IN2(n125), .IN3(N784), .IN4(n126), .IN5(N721), 
        .IN6(n127), .Q(n169) );
  AO222X1 U458 ( .IN1(N843), .IN2(n128), .IN3(N871), .IN4(n129), .IN5(N814), 
        .IN6(n130), .Q(n168) );
  AO222X1 U459 ( .IN1(N924), .IN2(n131), .IN3(N949), .IN4(n132), .IN5(N898), 
        .IN6(n133), .Q(n167) );
  AO222X1 U460 ( .IN1(N996), .IN2(n134), .IN3(N1018), .IN4(n135), .IN5(N973), 
        .IN6(n136), .Q(n166) );
  NOR4X0 U461 ( .IN1(n170), .IN2(n171), .IN3(n172), .IN4(n173), .QN(n164) );
  AO222X1 U462 ( .IN1(N302), .IN2(n141), .IN3(N345), .IN4(n142), .IN5(n84), 
        .IN6(add_sum[23]), .Q(n173) );
  AO222X1 U463 ( .IN1(N387), .IN2(n143), .IN3(N468), .IN4(n144), .IN5(N428), 
        .IN6(n145), .Q(n172) );
  AO222X1 U464 ( .IN1(N545), .IN2(n146), .IN3(N583), .IN4(n147), .IN5(N507), 
        .IN6(n148), .Q(n171) );
  AO222X1 U465 ( .IN1(N619), .IN2(n149), .IN3(N688), .IN4(n150), .IN5(N654), 
        .IN6(n151), .Q(n170) );
  AO222X1 U466 ( .IN1(N196), .IN2(n115), .IN3(n62), .IN4(n174), .IN5(n118), 
        .IN6(n80), .Q(add_updated_exponent[4]) );
  NAND2X0 U467 ( .IN1(n175), .IN2(n176), .QN(n174) );
  NOR4X0 U468 ( .IN1(n177), .IN2(n178), .IN3(n179), .IN4(n180), .QN(n176) );
  AO222X1 U469 ( .IN1(N752), .IN2(n125), .IN3(N783), .IN4(n126), .IN5(N720), 
        .IN6(n127), .Q(n180) );
  AO222X1 U470 ( .IN1(n81), .IN2(n128), .IN3(N870), .IN4(n129), .IN5(N813), 
        .IN6(n130), .Q(n179) );
  AO222X1 U471 ( .IN1(N923), .IN2(n131), .IN3(N948), .IN4(n132), .IN5(N897), 
        .IN6(n133), .Q(n178) );
  AO222X1 U472 ( .IN1(N995), .IN2(n134), .IN3(N1017), .IN4(n135), .IN5(N972), 
        .IN6(n136), .Q(n177) );
  NOR4X0 U473 ( .IN1(n181), .IN2(n182), .IN3(n183), .IN4(n184), .QN(n175) );
  AO222X1 U474 ( .IN1(N301), .IN2(n141), .IN3(N344), .IN4(n142), .IN5(
        add_sum[23]), .IN6(n80), .Q(n184) );
  AO222X1 U475 ( .IN1(N386), .IN2(n143), .IN3(N467), .IN4(n144), .IN5(N427), 
        .IN6(n145), .Q(n183) );
  AO222X1 U476 ( .IN1(N544), .IN2(n146), .IN3(N582), .IN4(n147), .IN5(N506), 
        .IN6(n148), .Q(n182) );
  AO222X1 U477 ( .IN1(N618), .IN2(n149), .IN3(N687), .IN4(n150), .IN5(N653), 
        .IN6(n151), .Q(n181) );
  AO222X1 U478 ( .IN1(N195), .IN2(n115), .IN3(n62), .IN4(n185), .IN5(n118), 
        .IN6(n75), .Q(add_updated_exponent[3]) );
  NAND2X0 U479 ( .IN1(n186), .IN2(n187), .QN(n185) );
  NOR4X0 U480 ( .IN1(n188), .IN2(n189), .IN3(n190), .IN4(n191), .QN(n187) );
  AO222X1 U481 ( .IN1(N751), .IN2(n125), .IN3(N782), .IN4(n126), .IN5(N719), 
        .IN6(n127), .Q(n191) );
  AO222X1 U482 ( .IN1(N922), .IN2(n131), .IN3(N947), .IN4(n132), .IN5(N896), 
        .IN6(n133), .Q(n189) );
  AO222X1 U483 ( .IN1(N994), .IN2(n134), .IN3(N1016), .IN4(n135), .IN5(N971), 
        .IN6(n136), .Q(n188) );
  NOR4X0 U484 ( .IN1(n192), .IN2(n193), .IN3(n194), .IN4(n195), .QN(n186) );
  AO222X1 U485 ( .IN1(N300), .IN2(n141), .IN3(N343), .IN4(n142), .IN5(
        add_sum[23]), .IN6(n76), .Q(n195) );
  AO222X1 U486 ( .IN1(N385), .IN2(n143), .IN3(N466), .IN4(n144), .IN5(N426), 
        .IN6(n145), .Q(n194) );
  AO222X1 U487 ( .IN1(N543), .IN2(n146), .IN3(n77), .IN4(n147), .IN5(N505), 
        .IN6(n148), .Q(n193) );
  AO222X1 U488 ( .IN1(N617), .IN2(n149), .IN3(N686), .IN4(n150), .IN5(N652), 
        .IN6(n151), .Q(n192) );
  AO222X1 U489 ( .IN1(N194), .IN2(n115), .IN3(n62), .IN4(n196), .IN5(n118), 
        .IN6(n73), .Q(add_updated_exponent[2]) );
  NAND2X0 U490 ( .IN1(n197), .IN2(n198), .QN(n196) );
  NOR4X0 U491 ( .IN1(n199), .IN2(n200), .IN3(n201), .IN4(n202), .QN(n198) );
  AO222X1 U492 ( .IN1(N750), .IN2(n125), .IN3(N781), .IN4(n126), .IN5(n74), 
        .IN6(n127), .Q(n202) );
  AO222X1 U493 ( .IN1(n73), .IN2(n128), .IN3(N868), .IN4(n129), .IN5(N811), 
        .IN6(n130), .Q(n201) );
  AO222X1 U494 ( .IN1(N921), .IN2(n131), .IN3(n74), .IN4(n132), .IN5(N895), 
        .IN6(n133), .Q(n200) );
  AO222X1 U495 ( .IN1(N993), .IN2(n134), .IN3(N1015), .IN4(n135), .IN5(N970), 
        .IN6(n136), .Q(n199) );
  NOR4X0 U496 ( .IN1(n203), .IN2(n204), .IN3(n205), .IN4(n206), .QN(n197) );
  AO222X1 U497 ( .IN1(N299), .IN2(n141), .IN3(N342), .IN4(n142), .IN5(
        add_sum[23]), .IN6(n73), .Q(n206) );
  AO222X1 U498 ( .IN1(N384), .IN2(n143), .IN3(N465), .IN4(n144), .IN5(n74), 
        .IN6(n145), .Q(n205) );
  AO222X1 U499 ( .IN1(N542), .IN2(n146), .IN3(n73), .IN4(n147), .IN5(N504), 
        .IN6(n148), .Q(n204) );
  AO222X1 U500 ( .IN1(N616), .IN2(n149), .IN3(N685), .IN4(n150), .IN5(N651), 
        .IN6(n151), .Q(n203) );
  AO222X1 U501 ( .IN1(N193), .IN2(n115), .IN3(n62), .IN4(n207), .IN5(n118), 
        .IN6(n69), .Q(add_updated_exponent[1]) );
  NAND2X0 U502 ( .IN1(n208), .IN2(n209), .QN(n207) );
  NOR4X0 U503 ( .IN1(n210), .IN2(n211), .IN3(n212), .IN4(n213), .QN(n209) );
  AO222X1 U504 ( .IN1(N749), .IN2(n125), .IN3(n70), .IN4(n126), .IN5(n69), 
        .IN6(n127), .Q(n213) );
  AO222X1 U505 ( .IN1(n69), .IN2(n128), .IN3(N867), .IN4(n129), .IN5(N810), 
        .IN6(n130), .Q(n212) );
  AO222X1 U506 ( .IN1(N920), .IN2(n131), .IN3(n69), .IN4(n132), .IN5(n70), 
        .IN6(n133), .Q(n211) );
  AO222X1 U507 ( .IN1(n70), .IN2(n134), .IN3(N1014), .IN4(n135), .IN5(N969), 
        .IN6(n136), .Q(n210) );
  NOR4X0 U508 ( .IN1(n214), .IN2(n215), .IN3(n216), .IN4(n217), .QN(n208) );
  AO222X1 U509 ( .IN1(N298), .IN2(n141), .IN3(n70), .IN4(n142), .IN5(
        add_sum[23]), .IN6(n69), .Q(n217) );
  AO222X1 U510 ( .IN1(N383), .IN2(n143), .IN3(N464), .IN4(n144), .IN5(N424), 
        .IN6(n145), .Q(n216) );
  AO222X1 U511 ( .IN1(N541), .IN2(n146), .IN3(n68), .IN4(n147), .IN5(n70), 
        .IN6(n148), .Q(n215) );
  AO222X1 U512 ( .IN1(N615), .IN2(n149), .IN3(N684), .IN4(n150), .IN5(n70), 
        .IN6(n151), .Q(n214) );
  AO222X1 U513 ( .IN1(N192), .IN2(n115), .IN3(n62), .IN4(n218), .IN5(n118), 
        .IN6(n65), .Q(add_updated_exponent[0]) );
  NAND2X0 U514 ( .IN1(n219), .IN2(n220), .QN(n218) );
  NOR4X0 U515 ( .IN1(n221), .IN2(n222), .IN3(n223), .IN4(n224), .QN(n220) );
  AO222X1 U516 ( .IN1(n67), .IN2(n125), .IN3(n65), .IN4(n126), .IN5(n65), 
        .IN6(n127), .Q(n224) );
  AO222X1 U517 ( .IN1(n66), .IN2(n128), .IN3(n67), .IN4(n129), .IN5(n67), 
        .IN6(n130), .Q(n223) );
  AO222X1 U518 ( .IN1(n67), .IN2(n131), .IN3(n65), .IN4(n132), .IN5(n65), 
        .IN6(n133), .Q(n222) );
  AO222X1 U519 ( .IN1(n66), .IN2(n134), .IN3(n67), .IN4(n135), .IN5(n67), 
        .IN6(n136), .Q(n221) );
  INVX0 U520 ( .INP(n225), .ZN(n135) );
  NOR4X0 U521 ( .IN1(n226), .IN2(n227), .IN3(n228), .IN4(n229), .QN(n219) );
  AO222X1 U522 ( .IN1(n67), .IN2(n141), .IN3(n65), .IN4(n142), .IN5(
        add_sum[23]), .IN6(n65), .Q(n229) );
  AO222X1 U523 ( .IN1(n67), .IN2(n143), .IN3(n67), .IN4(n144), .IN5(n65), 
        .IN6(n145), .Q(n228) );
  AO222X1 U524 ( .IN1(n67), .IN2(n146), .IN3(n65), .IN4(n147), .IN5(n65), 
        .IN6(n148), .Q(n227) );
  AO222X1 U525 ( .IN1(n67), .IN2(n149), .IN3(n67), .IN4(n150), .IN5(n65), 
        .IN6(n151), .Q(n226) );
  NAND2X0 U526 ( .IN1(n230), .IN2(n231), .QN(n115) );
  AO221X1 U527 ( .IN1(n62), .IN2(n232), .IN3(N210), .IN4(n233), .IN5(n234), 
        .Q(add_updated_add_sum[9]) );
  AO22X1 U528 ( .IN1(n235), .IN2(add_sum[10]), .IN3(n63), .IN4(add_sum[9]), 
        .Q(n234) );
  NAND4X0 U529 ( .IN1(n236), .IN2(n237), .IN3(n238), .IN4(n239), .QN(n232) );
  OA222X1 U530 ( .IN1(n240), .IN2(n241), .IN3(n242), .IN4(n243), .IN5(n244), 
        .IN6(n245), .Q(n239) );
  OA22X1 U531 ( .IN1(n246), .IN2(n247), .IN3(n248), .IN4(n249), .Q(n238) );
  OA222X1 U532 ( .IN1(n250), .IN2(n251), .IN3(n252), .IN4(n253), .IN5(n254), 
        .IN6(n255), .Q(n237) );
  OA22X1 U533 ( .IN1(n256), .IN2(n257), .IN3(n258), .IN4(n259), .Q(n236) );
  AO221X1 U534 ( .IN1(n116), .IN2(n260), .IN3(N209), .IN4(n64), .IN5(n261), 
        .Q(add_updated_add_sum[8]) );
  AO22X1 U535 ( .IN1(n235), .IN2(add_sum[9]), .IN3(n63), .IN4(add_sum[8]), .Q(
        n261) );
  NAND4X0 U536 ( .IN1(n262), .IN2(n263), .IN3(n264), .IN4(n265), .QN(n260) );
  AOI222X1 U537 ( .IN1(add_sum[2]), .IN2(n148), .IN3(n147), .IN4(add_sum[0]), 
        .IN5(add_sum[1]), .IN6(n146), .QN(n265) );
  OA22X1 U538 ( .IN1(n246), .IN2(n249), .IN3(n254), .IN4(n253), .Q(n264) );
  OA22X1 U539 ( .IN1(n248), .IN2(n255), .IN3(n252), .IN4(n251), .Q(n263) );
  OA22X1 U540 ( .IN1(n250), .IN2(n257), .IN3(n258), .IN4(n256), .Q(n262) );
  AO221X1 U541 ( .IN1(n116), .IN2(n266), .IN3(N208), .IN4(n64), .IN5(n267), 
        .Q(add_updated_add_sum[7]) );
  AO22X1 U542 ( .IN1(n235), .IN2(add_sum[8]), .IN3(n63), .IN4(add_sum[7]), .Q(
        n267) );
  NAND4X0 U543 ( .IN1(n268), .IN2(n269), .IN3(n270), .IN4(n271), .QN(n266) );
  OA22X1 U544 ( .IN1(n241), .IN2(n243), .IN3(n244), .IN4(n247), .Q(n271) );
  OA22X1 U545 ( .IN1(n240), .IN2(n249), .IN3(n248), .IN4(n253), .Q(n270) );
  OA22X1 U546 ( .IN1(n246), .IN2(n255), .IN3(n254), .IN4(n251), .Q(n269) );
  OA22X1 U547 ( .IN1(n252), .IN2(n257), .IN3(n258), .IN4(n250), .Q(n268) );
  AO221X1 U548 ( .IN1(n116), .IN2(n272), .IN3(N207), .IN4(n64), .IN5(n273), 
        .Q(add_updated_add_sum[6]) );
  AO22X1 U549 ( .IN1(n235), .IN2(add_sum[7]), .IN3(add_sum[6]), .IN4(n274), 
        .Q(n273) );
  NAND2X0 U550 ( .IN1(n275), .IN2(n276), .QN(n272) );
  AOI222X1 U551 ( .IN1(add_sum[3]), .IN2(n143), .IN3(n148), .IN4(add_sum[0]), 
        .IN5(add_sum[1]), .IN6(n144), .QN(n276) );
  AOI222X1 U552 ( .IN1(add_sum[5]), .IN2(n141), .IN3(add_sum[2]), .IN4(n145), 
        .IN5(add_sum[4]), .IN6(n142), .QN(n275) );
  AO221X1 U553 ( .IN1(n116), .IN2(n277), .IN3(N206), .IN4(n64), .IN5(n278), 
        .Q(add_updated_add_sum[5]) );
  AO22X1 U554 ( .IN1(n235), .IN2(add_sum[6]), .IN3(add_sum[5]), .IN4(n274), 
        .Q(n278) );
  AO221X1 U555 ( .IN1(n142), .IN2(add_sum[3]), .IN3(n141), .IN4(add_sum[4]), 
        .IN5(n279), .Q(n277) );
  AO222X1 U556 ( .IN1(n143), .IN2(add_sum[2]), .IN3(add_sum[0]), .IN4(n144), 
        .IN5(n145), .IN6(add_sum[1]), .Q(n279) );
  AO221X1 U557 ( .IN1(n116), .IN2(n280), .IN3(N205), .IN4(n64), .IN5(n281), 
        .Q(add_updated_add_sum[4]) );
  AO22X1 U558 ( .IN1(n235), .IN2(add_sum[5]), .IN3(add_sum[4]), .IN4(n274), 
        .Q(n281) );
  AO221X1 U559 ( .IN1(n142), .IN2(add_sum[2]), .IN3(n141), .IN4(add_sum[3]), 
        .IN5(n282), .Q(n280) );
  AO22X1 U560 ( .IN1(add_sum[0]), .IN2(n145), .IN3(n143), .IN4(add_sum[1]), 
        .Q(n282) );
  AO221X1 U561 ( .IN1(n116), .IN2(n283), .IN3(N204), .IN4(n64), .IN5(n284), 
        .Q(add_updated_add_sum[3]) );
  AO22X1 U562 ( .IN1(n235), .IN2(add_sum[4]), .IN3(add_sum[3]), .IN4(n274), 
        .Q(n284) );
  AO222X1 U563 ( .IN1(n142), .IN2(add_sum[1]), .IN3(add_sum[0]), .IN4(n143), 
        .IN5(n141), .IN6(add_sum[2]), .Q(n283) );
  AO221X1 U564 ( .IN1(n116), .IN2(n285), .IN3(N203), .IN4(n64), .IN5(n286), 
        .Q(add_updated_add_sum[2]) );
  AO22X1 U565 ( .IN1(n235), .IN2(add_sum[3]), .IN3(add_sum[2]), .IN4(n274), 
        .Q(n286) );
  AO22X1 U566 ( .IN1(n141), .IN2(add_sum[1]), .IN3(add_sum[0]), .IN4(n142), 
        .Q(n285) );
  AND2X1 U567 ( .IN1(N225), .IN2(n64), .Q(add_updated_add_sum[24]) );
  AO221X1 U568 ( .IN1(N224), .IN2(n64), .IN3(add_sum[24]), .IN4(n235), .IN5(
        n287), .Q(add_updated_add_sum[23]) );
  AO21X1 U569 ( .IN1(n62), .IN2(n288), .IN3(n118), .Q(n287) );
  NAND4X0 U570 ( .IN1(n289), .IN2(n290), .IN3(n291), .IN4(n292), .QN(n288) );
  NOR4X0 U571 ( .IN1(n293), .IN2(n134), .IN3(add_sum[23]), .IN4(n136), .QN(
        n292) );
  NAND3X0 U572 ( .IN1(n257), .IN2(n225), .IN3(n251), .QN(n293) );
  NAND3X0 U573 ( .IN1(n294), .IN2(n295), .IN3(n296), .QN(n225) );
  NOR4X0 U574 ( .IN1(n297), .IN2(n144), .IN3(n145), .IN4(n143), .QN(n291) );
  NAND3X0 U575 ( .IN1(n241), .IN2(n247), .IN3(n245), .QN(n297) );
  NOR4X0 U576 ( .IN1(n298), .IN2(n126), .IN3(n127), .IN4(n125), .QN(n290) );
  NAND3X0 U577 ( .IN1(n242), .IN2(n299), .IN3(n300), .QN(n298) );
  NOR4X0 U578 ( .IN1(n301), .IN2(n129), .IN3(n130), .IN4(n128), .QN(n289) );
  NAND3X0 U579 ( .IN1(n302), .IN2(n303), .IN3(n304), .QN(n301) );
  AO221X1 U580 ( .IN1(n116), .IN2(n305), .IN3(N223), .IN4(n64), .IN5(n306), 
        .Q(add_updated_add_sum[22]) );
  AO22X1 U581 ( .IN1(n235), .IN2(add_sum[23]), .IN3(n63), .IN4(add_sum[22]), 
        .Q(n306) );
  NAND4X0 U582 ( .IN1(n307), .IN2(n308), .IN3(n309), .IN4(n310), .QN(n305) );
  NOR4X0 U583 ( .IN1(n311), .IN2(n312), .IN3(n313), .IN4(n314), .QN(n310) );
  AO222X1 U584 ( .IN1(n127), .IN2(add_sum[10]), .IN3(n125), .IN4(add_sum[9]), 
        .IN5(n150), .IN6(add_sum[11]), .Q(n314) );
  AO222X1 U585 ( .IN1(n130), .IN2(add_sum[7]), .IN3(n128), .IN4(add_sum[6]), 
        .IN5(n126), .IN6(add_sum[8]), .Q(n313) );
  INVX0 U586 ( .INP(n315), .ZN(n128) );
  INVX0 U587 ( .INP(n316), .ZN(n130) );
  AO222X1 U588 ( .IN1(n133), .IN2(add_sum[4]), .IN3(n131), .IN4(add_sum[3]), 
        .IN5(n129), .IN6(add_sum[5]), .Q(n312) );
  INVX0 U589 ( .INP(n317), .ZN(n129) );
  INVX0 U590 ( .INP(n302), .ZN(n131) );
  INVX0 U591 ( .INP(n303), .ZN(n133) );
  AO222X1 U592 ( .IN1(n136), .IN2(add_sum[1]), .IN3(add_sum[0]), .IN4(n134), 
        .IN5(n132), .IN6(add_sum[2]), .Q(n311) );
  INVX0 U593 ( .INP(n304), .ZN(n132) );
  INVX0 U594 ( .INP(n319), .ZN(n136) );
  OA221X1 U595 ( .IN1(n258), .IN2(n320), .IN3(n321), .IN4(n257), .IN5(n322), 
        .Q(n309) );
  OA222X1 U596 ( .IN1(n323), .IN2(n251), .IN3(n253), .IN4(n324), .IN5(n325), 
        .IN6(n255), .Q(n322) );
  OA222X1 U597 ( .IN1(n326), .IN2(n245), .IN3(n242), .IN4(n327), .IN5(n328), 
        .IN6(n299), .Q(n308) );
  OA222X1 U598 ( .IN1(n329), .IN2(n249), .IN3(n330), .IN4(n241), .IN5(n331), 
        .IN6(n247), .Q(n307) );
  AO221X1 U599 ( .IN1(n116), .IN2(n332), .IN3(N222), .IN4(n64), .IN5(n333), 
        .Q(add_updated_add_sum[21]) );
  AO22X1 U600 ( .IN1(n235), .IN2(add_sum[22]), .IN3(n63), .IN4(add_sum[21]), 
        .Q(n333) );
  NAND4X0 U601 ( .IN1(n334), .IN2(n335), .IN3(n336), .IN4(n337), .QN(n332) );
  AND4X1 U602 ( .IN1(n338), .IN2(n339), .IN3(n340), .IN4(n341), .Q(n337) );
  AOI222X1 U603 ( .IN1(add_sum[13]), .IN2(n147), .IN3(add_sum[12]), .IN4(n149), 
        .IN5(add_sum[11]), .IN6(n151), .QN(n341) );
  INVX0 U604 ( .INP(n242), .ZN(n149) );
  OA222X1 U605 ( .IN1(n331), .IN2(n249), .IN3(n326), .IN4(n241), .IN5(n330), 
        .IN6(n247), .Q(n340) );
  OA222X1 U606 ( .IN1(n324), .IN2(n251), .IN3(n325), .IN4(n253), .IN5(n329), 
        .IN6(n255), .Q(n339) );
  OA22X1 U607 ( .IN1(n323), .IN2(n257), .IN3(n258), .IN4(n321), .Q(n338) );
  OA221X1 U608 ( .IN1(n342), .IN2(n300), .IN3(n259), .IN4(n343), .IN5(n344), 
        .Q(n336) );
  OA222X1 U609 ( .IN1(n256), .IN2(n345), .IN3(n252), .IN4(n316), .IN5(n250), 
        .IN6(n346), .Q(n344) );
  OA222X1 U610 ( .IN1(n240), .IN2(n302), .IN3(n319), .IN4(n243), .IN5(n244), 
        .IN6(n304), .Q(n335) );
  NAND3X0 U611 ( .IN1(n296), .IN2(n318), .IN3(add_sum[2]), .QN(n319) );
  OA222X1 U612 ( .IN1(n254), .IN2(n315), .IN3(n246), .IN4(n303), .IN5(n248), 
        .IN6(n317), .Q(n334) );
  AO221X1 U613 ( .IN1(n116), .IN2(n347), .IN3(N221), .IN4(n64), .IN5(n348), 
        .Q(add_updated_add_sum[20]) );
  AO22X1 U614 ( .IN1(n235), .IN2(add_sum[21]), .IN3(n63), .IN4(add_sum[20]), 
        .Q(n348) );
  NAND4X0 U615 ( .IN1(n349), .IN2(n350), .IN3(n351), .IN4(n352), .QN(n347) );
  NOR2X0 U616 ( .IN1(n353), .IN2(n354), .QN(n352) );
  AO221X1 U617 ( .IN1(n141), .IN2(add_sum[19]), .IN3(add_sum[20]), .IN4(n355), 
        .IN5(n356), .Q(n354) );
  AO222X1 U618 ( .IN1(n145), .IN2(add_sum[16]), .IN3(n143), .IN4(add_sum[17]), 
        .IN5(n142), .IN6(add_sum[18]), .Q(n356) );
  AO221X1 U619 ( .IN1(n148), .IN2(add_sum[14]), .IN3(n144), .IN4(add_sum[15]), 
        .IN5(n357), .Q(n353) );
  AO222X1 U620 ( .IN1(n147), .IN2(add_sum[12]), .IN3(n151), .IN4(add_sum[10]), 
        .IN5(n146), .IN6(add_sum[13]), .Q(n357) );
  OA221X1 U621 ( .IN1(n358), .IN2(n242), .IN3(n259), .IN4(n300), .IN5(n359), 
        .Q(n351) );
  AOI222X1 U622 ( .IN1(add_sum[8]), .IN2(n127), .IN3(add_sum[6]), .IN4(n126), 
        .IN5(add_sum[7]), .IN6(n125), .QN(n359) );
  INVX0 U623 ( .INP(n346), .ZN(n126) );
  OA222X1 U624 ( .IN1(n240), .IN2(n303), .IN3(n304), .IN4(n243), .IN5(n244), 
        .IN6(n302), .Q(n350) );
  NAND4X0 U625 ( .IN1(add_sum[3]), .IN2(n360), .IN3(n361), .IN4(n362), .QN(
        n304) );
  INVX0 U626 ( .INP(n363), .ZN(n362) );
  OA222X1 U627 ( .IN1(n254), .IN2(n316), .IN3(n246), .IN4(n317), .IN5(n248), 
        .IN6(n315), .Q(n349) );
  AO221X1 U628 ( .IN1(n364), .IN2(add_sum[0]), .IN3(N202), .IN4(n64), .IN5(
        n365), .Q(add_updated_add_sum[1]) );
  AO22X1 U629 ( .IN1(n235), .IN2(add_sum[2]), .IN3(add_sum[1]), .IN4(n274), 
        .Q(n365) );
  NOR2X0 U630 ( .IN1(n366), .IN2(n257), .QN(n364) );
  AO221X1 U631 ( .IN1(n116), .IN2(n367), .IN3(N220), .IN4(n233), .IN5(n368), 
        .Q(add_updated_add_sum[19]) );
  AO22X1 U632 ( .IN1(n235), .IN2(add_sum[20]), .IN3(n63), .IN4(add_sum[19]), 
        .Q(n368) );
  NAND4X0 U633 ( .IN1(n369), .IN2(n370), .IN3(n371), .IN4(n372), .QN(n367) );
  OA221X1 U634 ( .IN1(n248), .IN2(n316), .IN3(n246), .IN4(n315), .IN5(n373), 
        .Q(n372) );
  OA222X1 U635 ( .IN1(n240), .IN2(n317), .IN3(n302), .IN4(n243), .IN5(n244), 
        .IN6(n303), .Q(n373) );
  NAND4X0 U636 ( .IN1(add_sum[4]), .IN2(n360), .IN3(n374), .IN4(n254), .QN(
        n302) );
  OA221X1 U637 ( .IN1(n342), .IN2(n242), .IN3(n256), .IN4(n300), .IN5(n375), 
        .Q(n371) );
  OA222X1 U638 ( .IN1(n250), .IN2(n343), .IN3(n254), .IN4(n346), .IN5(n252), 
        .IN6(n345), .Q(n375) );
  OA221X1 U639 ( .IN1(n326), .IN2(n249), .IN3(n327), .IN4(n247), .IN5(n376), 
        .Q(n370) );
  OA222X1 U640 ( .IN1(n328), .IN2(n241), .IN3(n259), .IN4(n299), .IN5(n358), 
        .IN6(n245), .Q(n376) );
  OA221X1 U641 ( .IN1(n258), .IN2(n324), .IN3(n325), .IN4(n257), .IN5(n377), 
        .Q(n369) );
  OA222X1 U642 ( .IN1(n329), .IN2(n251), .IN3(n331), .IN4(n253), .IN5(n330), 
        .IN6(n255), .Q(n377) );
  AO221X1 U643 ( .IN1(n116), .IN2(n378), .IN3(N219), .IN4(n233), .IN5(n379), 
        .Q(add_updated_add_sum[18]) );
  AO22X1 U644 ( .IN1(n235), .IN2(add_sum[19]), .IN3(n63), .IN4(add_sum[18]), 
        .Q(n379) );
  NAND4X0 U645 ( .IN1(n380), .IN2(n381), .IN3(n382), .IN4(n383), .QN(n378) );
  OA221X1 U646 ( .IN1(n248), .IN2(n346), .IN3(n246), .IN4(n316), .IN5(n384), 
        .Q(n383) );
  OA222X1 U647 ( .IN1(n240), .IN2(n315), .IN3(n303), .IN4(n243), .IN5(n244), 
        .IN6(n317), .Q(n384) );
  NAND3X0 U648 ( .IN1(n360), .IN2(n385), .IN3(add_sum[5]), .QN(n303) );
  INVX0 U649 ( .INP(n386), .ZN(n385) );
  OA221X1 U650 ( .IN1(n256), .IN2(n299), .IN3(n259), .IN4(n242), .IN5(n387), 
        .Q(n382) );
  AOI222X1 U651 ( .IN1(add_sum[7]), .IN2(n150), .IN3(add_sum[5]), .IN4(n125), 
        .IN5(add_sum[6]), .IN6(n127), .QN(n387) );
  INVX0 U652 ( .INP(n343), .ZN(n127) );
  INVX0 U653 ( .INP(n345), .ZN(n125) );
  INVX0 U654 ( .INP(n300), .ZN(n150) );
  OA221X1 U655 ( .IN1(n330), .IN2(n253), .IN3(n327), .IN4(n249), .IN5(n388), 
        .Q(n381) );
  OA222X1 U656 ( .IN1(n328), .IN2(n247), .IN3(n342), .IN4(n245), .IN5(n358), 
        .IN6(n241), .Q(n388) );
  OA221X1 U657 ( .IN1(n331), .IN2(n251), .IN3(n326), .IN4(n255), .IN5(n389), 
        .Q(n380) );
  OA22X1 U658 ( .IN1(n329), .IN2(n257), .IN3(n258), .IN4(n325), .Q(n389) );
  AO221X1 U659 ( .IN1(n116), .IN2(n390), .IN3(N218), .IN4(n233), .IN5(n391), 
        .Q(add_updated_add_sum[17]) );
  AO22X1 U660 ( .IN1(n235), .IN2(add_sum[18]), .IN3(n63), .IN4(add_sum[17]), 
        .Q(n391) );
  NAND4X0 U661 ( .IN1(n392), .IN2(n393), .IN3(n394), .IN4(n395), .QN(n390) );
  OA221X1 U662 ( .IN1(n248), .IN2(n345), .IN3(n246), .IN4(n346), .IN5(n396), 
        .Q(n395) );
  OA222X1 U663 ( .IN1(n240), .IN2(n316), .IN3(n317), .IN4(n243), .IN5(n244), 
        .IN6(n315), .Q(n396) );
  NAND3X0 U664 ( .IN1(n397), .IN2(n398), .IN3(add_sum[6]), .QN(n317) );
  INVX0 U665 ( .INP(n399), .ZN(n398) );
  OA221X1 U666 ( .IN1(n252), .IN2(n300), .IN3(n254), .IN4(n343), .IN5(n400), 
        .Q(n394) );
  OA22X1 U667 ( .IN1(n256), .IN2(n242), .IN3(n250), .IN4(n299), .Q(n400) );
  OA221X1 U668 ( .IN1(n326), .IN2(n253), .IN3(n328), .IN4(n249), .IN5(n401), 
        .Q(n393) );
  AOI222X1 U669 ( .IN1(add_sum[11]), .IN2(n148), .IN3(add_sum[9]), .IN4(n147), 
        .IN5(add_sum[10]), .IN6(n146), .QN(n401) );
  OA221X1 U670 ( .IN1(n330), .IN2(n251), .IN3(n327), .IN4(n255), .IN5(n402), 
        .Q(n392) );
  OA22X1 U671 ( .IN1(n331), .IN2(n257), .IN3(n258), .IN4(n329), .Q(n402) );
  AO221X1 U672 ( .IN1(n116), .IN2(n403), .IN3(N217), .IN4(n233), .IN5(n404), 
        .Q(add_updated_add_sum[16]) );
  AO22X1 U673 ( .IN1(n235), .IN2(add_sum[17]), .IN3(n63), .IN4(add_sum[16]), 
        .Q(n404) );
  NAND4X0 U674 ( .IN1(n405), .IN2(n406), .IN3(n407), .IN4(n408), .QN(n403) );
  OA221X1 U675 ( .IN1(n248), .IN2(n343), .IN3(n246), .IN4(n345), .IN5(n409), 
        .Q(n408) );
  OA222X1 U676 ( .IN1(n240), .IN2(n346), .IN3(n315), .IN4(n243), .IN5(n244), 
        .IN6(n316), .Q(n409) );
  NAND4X0 U677 ( .IN1(add_sum[7]), .IN2(n410), .IN3(n411), .IN4(n412), .QN(
        n315) );
  NOR2X0 U678 ( .IN1(add_sum[9]), .IN2(add_sum[8]), .QN(n411) );
  OA221X1 U679 ( .IN1(n256), .IN2(n245), .IN3(n252), .IN4(n299), .IN5(n413), 
        .Q(n407) );
  OA22X1 U680 ( .IN1(n254), .IN2(n300), .IN3(n250), .IN4(n242), .Q(n413) );
  OA221X1 U681 ( .IN1(n342), .IN2(n247), .IN3(n259), .IN4(n241), .IN5(n414), 
        .Q(n406) );
  OA22X1 U682 ( .IN1(n358), .IN2(n249), .IN3(n327), .IN4(n253), .Q(n414) );
  OA221X1 U683 ( .IN1(n326), .IN2(n251), .IN3(n328), .IN4(n255), .IN5(n415), 
        .Q(n405) );
  OA22X1 U684 ( .IN1(n330), .IN2(n257), .IN3(n258), .IN4(n331), .Q(n415) );
  AO221X1 U685 ( .IN1(n116), .IN2(n416), .IN3(N216), .IN4(n64), .IN5(n417), 
        .Q(add_updated_add_sum[15]) );
  AO22X1 U686 ( .IN1(n235), .IN2(add_sum[16]), .IN3(n63), .IN4(add_sum[15]), 
        .Q(n417) );
  NAND4X0 U687 ( .IN1(n418), .IN2(n419), .IN3(n420), .IN4(n421), .QN(n416) );
  OA221X1 U688 ( .IN1(n244), .IN2(n346), .IN3(n316), .IN4(n243), .IN5(n422), 
        .Q(n421) );
  OA22X1 U689 ( .IN1(n240), .IN2(n345), .IN3(n246), .IN4(n343), .Q(n422) );
  NAND4X0 U690 ( .IN1(add_sum[8]), .IN2(n410), .IN3(n423), .IN4(n259), .QN(
        n316) );
  INVX0 U691 ( .INP(n424), .ZN(n423) );
  OA221X1 U692 ( .IN1(n250), .IN2(n245), .IN3(n254), .IN4(n299), .IN5(n425), 
        .Q(n420) );
  OA22X1 U693 ( .IN1(n248), .IN2(n300), .IN3(n252), .IN4(n242), .Q(n425) );
  OA221X1 U694 ( .IN1(n259), .IN2(n247), .IN3(n256), .IN4(n241), .IN5(n426), 
        .Q(n419) );
  OA22X1 U695 ( .IN1(n342), .IN2(n249), .IN3(n328), .IN4(n253), .Q(n426) );
  OA221X1 U696 ( .IN1(n327), .IN2(n251), .IN3(n358), .IN4(n255), .IN5(n427), 
        .Q(n418) );
  OA22X1 U697 ( .IN1(n326), .IN2(n257), .IN3(n258), .IN4(n330), .Q(n427) );
  AO221X1 U698 ( .IN1(n116), .IN2(n428), .IN3(N215), .IN4(n233), .IN5(n429), 
        .Q(add_updated_add_sum[14]) );
  AO22X1 U699 ( .IN1(n235), .IN2(add_sum[15]), .IN3(n63), .IN4(add_sum[14]), 
        .Q(n429) );
  NAND4X0 U700 ( .IN1(n430), .IN2(n431), .IN3(n432), .IN4(n433), .QN(n428) );
  OA221X1 U701 ( .IN1(n244), .IN2(n345), .IN3(n346), .IN4(n243), .IN5(n434), 
        .Q(n433) );
  OA22X1 U702 ( .IN1(n240), .IN2(n343), .IN3(n246), .IN4(n300), .Q(n434) );
  NAND3X0 U703 ( .IN1(n410), .IN2(n435), .IN3(add_sum[9]), .QN(n346) );
  INVX0 U704 ( .INP(n436), .ZN(n435) );
  OA221X1 U705 ( .IN1(n248), .IN2(n299), .IN3(n254), .IN4(n242), .IN5(n437), 
        .Q(n432) );
  OA22X1 U706 ( .IN1(n252), .IN2(n245), .IN3(n250), .IN4(n241), .Q(n437) );
  OA221X1 U707 ( .IN1(n259), .IN2(n249), .IN3(n256), .IN4(n247), .IN5(n438), 
        .Q(n431) );
  OA22X1 U708 ( .IN1(n358), .IN2(n253), .IN3(n342), .IN4(n255), .Q(n438) );
  OA222X1 U709 ( .IN1(n258), .IN2(n326), .IN3(n328), .IN4(n251), .IN5(n327), 
        .IN6(n257), .Q(n430) );
  AO221X1 U710 ( .IN1(n116), .IN2(n439), .IN3(N214), .IN4(n233), .IN5(n440), 
        .Q(add_updated_add_sum[13]) );
  AO22X1 U711 ( .IN1(n235), .IN2(add_sum[14]), .IN3(n63), .IN4(add_sum[13]), 
        .Q(n440) );
  NAND4X0 U712 ( .IN1(n441), .IN2(n442), .IN3(n443), .IN4(n444), .QN(n439) );
  OA221X1 U713 ( .IN1(n244), .IN2(n343), .IN3(n345), .IN4(n243), .IN5(n445), 
        .Q(n444) );
  OA22X1 U714 ( .IN1(n240), .IN2(n300), .IN3(n248), .IN4(n242), .Q(n445) );
  NAND4X0 U715 ( .IN1(add_sum[10]), .IN2(n446), .IN3(n447), .IN4(n358), .QN(
        n345) );
  INVX0 U716 ( .INP(n448), .ZN(n447) );
  AOI222X1 U717 ( .IN1(add_sum[6]), .IN2(n146), .IN3(add_sum[3]), .IN4(n151), 
        .IN5(add_sum[5]), .IN6(n147), .QN(n443) );
  INVX0 U718 ( .INP(n245), .ZN(n147) );
  INVX0 U719 ( .INP(n299), .ZN(n151) );
  OA221X1 U720 ( .IN1(n256), .IN2(n249), .IN3(n250), .IN4(n247), .IN5(n449), 
        .Q(n442) );
  OA22X1 U721 ( .IN1(n342), .IN2(n253), .IN3(n259), .IN4(n255), .Q(n449) );
  OA222X1 U722 ( .IN1(n258), .IN2(n327), .IN3(n358), .IN4(n251), .IN5(n328), 
        .IN6(n257), .Q(n441) );
  INVX0 U723 ( .INP(add_sum[13]), .ZN(n327) );
  AO221X1 U724 ( .IN1(n62), .IN2(n450), .IN3(N213), .IN4(n233), .IN5(n451), 
        .Q(add_updated_add_sum[12]) );
  AO22X1 U725 ( .IN1(n235), .IN2(add_sum[13]), .IN3(n63), .IN4(add_sum[12]), 
        .Q(n451) );
  NAND4X0 U726 ( .IN1(n452), .IN2(n453), .IN3(n454), .IN4(n455), .QN(n450) );
  OA221X1 U727 ( .IN1(n244), .IN2(n300), .IN3(n343), .IN4(n243), .IN5(n456), 
        .Q(n455) );
  OA22X1 U728 ( .IN1(n246), .IN2(n242), .IN3(n240), .IN4(n299), .Q(n456) );
  OA222X1 U729 ( .IN1(n252), .IN2(n247), .IN3(n248), .IN4(n245), .IN5(n254), 
        .IN6(n241), .Q(n454) );
  AOI222X1 U730 ( .IN1(add_sum[8]), .IN2(n145), .IN3(add_sum[7]), .IN4(n144), 
        .IN5(add_sum[9]), .IN6(n143), .QN(n453) );
  INVX0 U731 ( .INP(n253), .ZN(n143) );
  INVX0 U732 ( .INP(n255), .ZN(n145) );
  OA222X1 U733 ( .IN1(n258), .IN2(n328), .IN3(n342), .IN4(n251), .IN5(n358), 
        .IN6(n257), .Q(n452) );
  AO221X1 U734 ( .IN1(n62), .IN2(n458), .IN3(N212), .IN4(n233), .IN5(n459), 
        .Q(add_updated_add_sum[11]) );
  AO22X1 U735 ( .IN1(n235), .IN2(add_sum[12]), .IN3(n118), .IN4(add_sum[11]), 
        .Q(n459) );
  NAND4X0 U736 ( .IN1(n460), .IN2(n461), .IN3(n462), .IN4(n463), .QN(n458) );
  OA222X1 U737 ( .IN1(n244), .IN2(n299), .IN3(n300), .IN4(n243), .IN5(n240), 
        .IN6(n242), .Q(n463) );
  NAND4X0 U738 ( .IN1(add_sum[12]), .IN2(n464), .IN3(n465), .IN4(n466), .QN(
        n300) );
  INVX0 U739 ( .INP(n467), .ZN(n466) );
  OA222X1 U740 ( .IN1(n254), .IN2(n247), .IN3(n246), .IN4(n245), .IN5(n248), 
        .IN6(n241), .Q(n462) );
  INVX0 U741 ( .INP(add_sum[4]), .ZN(n248) );
  OA222X1 U742 ( .IN1(n250), .IN2(n255), .IN3(n252), .IN4(n249), .IN5(n256), 
        .IN6(n253), .Q(n461) );
  AOI222X1 U743 ( .IN1(n355), .IN2(add_sum[11]), .IN3(add_sum[9]), .IN4(n142), 
        .IN5(add_sum[10]), .IN6(n141), .QN(n460) );
  AO221X1 U744 ( .IN1(n62), .IN2(n468), .IN3(N211), .IN4(n233), .IN5(n469), 
        .Q(add_updated_add_sum[10]) );
  AO22X1 U745 ( .IN1(n235), .IN2(add_sum[11]), .IN3(n118), .IN4(add_sum[10]), 
        .Q(n469) );
  NAND4X0 U746 ( .IN1(n470), .IN2(n471), .IN3(n472), .IN4(n473), .QN(n468) );
  OA222X1 U747 ( .IN1(n240), .IN2(n245), .IN3(n244), .IN4(n242), .IN5(n299), 
        .IN6(n243), .Q(n473) );
  NAND4X0 U748 ( .IN1(add_sum[13]), .IN2(n464), .IN3(n474), .IN4(n326), .QN(
        n299) );
  INVX0 U749 ( .INP(n476), .ZN(n475) );
  INVX0 U750 ( .INP(add_sum[1]), .ZN(n244) );
  NAND2X0 U751 ( .IN1(n479), .IN2(n77), .QN(n478) );
  INVX0 U752 ( .INP(add_sum[2]), .ZN(n240) );
  AOI222X1 U753 ( .IN1(add_sum[5]), .IN2(n144), .IN3(add_sum[3]), .IN4(n146), 
        .IN5(add_sum[4]), .IN6(n148), .QN(n472) );
  INVX0 U754 ( .INP(n247), .ZN(n148) );
  NAND4X0 U755 ( .IN1(add_sum[17]), .IN2(n480), .IN3(n481), .IN4(n325), .QN(
        n247) );
  INVX0 U756 ( .INP(n241), .ZN(n146) );
  NAND4X0 U757 ( .IN1(add_sum[16]), .IN2(n480), .IN3(n482), .IN4(n483), .QN(
        n241) );
  INVX0 U758 ( .INP(n249), .ZN(n144) );
  OA222X1 U759 ( .IN1(n256), .IN2(n251), .IN3(n250), .IN4(n253), .IN5(n252), 
        .IN6(n255), .Q(n471) );
  NAND2X0 U760 ( .IN1(n487), .IN2(n479), .QN(n486) );
  NAND4X0 U761 ( .IN1(add_sum[20]), .IN2(n258), .IN3(n488), .IN4(n489), .QN(
        n253) );
  NOR2X0 U762 ( .IN1(add_sum[22]), .IN2(add_sum[21]), .QN(n488) );
  INVX0 U763 ( .INP(n142), .ZN(n251) );
  OA22X1 U764 ( .IN1(n259), .IN2(n257), .IN3(n258), .IN4(n342), .Q(n470) );
  INVX0 U765 ( .INP(n355), .ZN(n258) );
  INVX0 U766 ( .INP(n141), .ZN(n257) );
  NOR3X0 U767 ( .IN1(n355), .IN2(n491), .IN3(n320), .QN(n141) );
  AO222X1 U768 ( .IN1(add_sum[0]), .IN2(n274), .IN3(N201), .IN4(n64), .IN5(
        n235), .IN6(add_sum[1]), .Q(add_updated_add_sum[0]) );
  INVX0 U769 ( .INP(n230), .ZN(n235) );
  NAND2X0 U770 ( .IN1(n492), .IN2(n243), .QN(n230) );
  INVX0 U771 ( .INP(add_sum[0]), .ZN(n243) );
  INVX0 U772 ( .INP(n231), .ZN(n233) );
  NAND2X0 U773 ( .IN1(add_sum[0]), .IN2(n492), .QN(n231) );
  AOI21X1 U774 ( .IN1(add_sum[23]), .IN2(n493), .IN3(n62), .QN(n492) );
  AO21X1 U775 ( .IN1(n62), .IN2(n355), .IN3(n118), .Q(n274) );
  AND3X1 U776 ( .IN1(add_sum[23]), .IN2(n493), .IN3(n366), .Q(n118) );
  INVX0 U777 ( .INP(add_sum[24]), .ZN(n493) );
  OA21X1 U778 ( .IN1(n494), .IN2(n495), .IN3(n116), .Q(add_exception2) );
  INVX0 U779 ( .INP(n366), .ZN(n116) );
  AO221X1 U780 ( .IN1(n496), .IN2(n497), .IN3(n360), .IN4(n498), .IN5(n499), 
        .Q(n495) );
  AO22X1 U781 ( .IN1(n480), .IN2(n500), .IN3(n464), .IN4(n501), .Q(n499) );
  AO221X1 U782 ( .IN1(n467), .IN2(n465), .IN3(n502), .IN4(n326), .IN5(n476), 
        .Q(n501) );
  OA21X1 U783 ( .IN1(n77), .IN2(n67), .IN3(n502), .Q(n476) );
  INVX0 U784 ( .INP(add_sum[14]), .ZN(n326) );
  INVX0 U785 ( .INP(n474), .ZN(n502) );
  NAND2X0 U786 ( .IN1(n503), .IN2(n504), .QN(n474) );
  OA21X1 U787 ( .IN1(n504), .IN2(n67), .IN3(n503), .Q(n467) );
  OAI221X1 U788 ( .IN1(n483), .IN2(n505), .IN3(n481), .IN4(add_sum[18]), .IN5(
        n484), .QN(n500) );
  OR2X1 U789 ( .IN1(n481), .IN2(n506), .Q(n484) );
  NAND2X0 U790 ( .IN1(n507), .IN2(n479), .QN(n481) );
  NAND3X0 U791 ( .IN1(n508), .IN2(n77), .IN3(n479), .QN(n483) );
  NAND2X0 U792 ( .IN1(n506), .IN2(n69), .QN(n508) );
  AO221X1 U793 ( .IN1(n363), .IN2(n361), .IN3(n509), .IN4(n254), .IN5(n386), 
        .Q(n498) );
  INVX0 U794 ( .INP(add_sum[5]), .ZN(n254) );
  INVX0 U795 ( .INP(n374), .ZN(n509) );
  NAND2X0 U796 ( .IN1(n363), .IN2(n510), .QN(n374) );
  NAND3X0 U797 ( .IN1(n80), .IN2(N424), .IN3(n65), .QN(n510) );
  OA22X1 U798 ( .IN1(n490), .IN2(n321), .IN3(n491), .IN4(n320), .Q(n497) );
  NOR2X0 U799 ( .IN1(n355), .IN2(n489), .QN(n496) );
  NAND3X0 U800 ( .IN1(n479), .IN2(n511), .IN3(n487), .QN(n489) );
  NAND2X0 U801 ( .IN1(n66), .IN2(n69), .QN(n511) );
  NAND4X0 U802 ( .IN1(n512), .IN2(n513), .IN3(n514), .IN4(n515), .QN(n494) );
  NAND3X0 U803 ( .IN1(n516), .IN2(n77), .IN3(n479), .QN(n515) );
  AO21X1 U804 ( .IN1(n485), .IN2(n74), .IN3(n477), .Q(n516) );
  NAND2X0 U805 ( .IN1(n399), .IN2(n397), .QN(n514) );
  OA21X1 U806 ( .IN1(n67), .IN2(n81), .IN3(n386), .Q(n399) );
  OA21X1 U807 ( .IN1(n81), .IN2(n70), .IN3(n363), .Q(n386) );
  OA21X1 U808 ( .IN1(n81), .IN2(n487), .IN3(n517), .Q(n363) );
  NAND3X0 U809 ( .IN1(n296), .IN2(n518), .IN3(n519), .QN(n513) );
  NAND2X0 U810 ( .IN1(n318), .IN2(n520), .QN(n518) );
  INVX0 U811 ( .INP(n294), .ZN(n520) );
  AO21X1 U812 ( .IN1(n506), .IN2(n80), .IN3(n295), .Q(n318) );
  INVX0 U813 ( .INP(n519), .ZN(n295) );
  OA21X1 U814 ( .IN1(n81), .IN2(n507), .IN3(n517), .Q(n519) );
  OA21X1 U815 ( .IN1(n74), .IN2(n70), .IN3(n77), .Q(n507) );
  AND3X1 U816 ( .IN1(n361), .IN2(n246), .IN3(n360), .Q(n296) );
  AND2X1 U817 ( .IN1(n397), .IN2(n252), .Q(n360) );
  INVX0 U818 ( .INP(add_sum[6]), .ZN(n252) );
  AND4X1 U819 ( .IN1(n410), .IN2(n250), .IN3(n256), .IN4(n259), .Q(n397) );
  AND3X1 U820 ( .IN1(n342), .IN2(n358), .IN3(n446), .Q(n410) );
  INVX0 U821 ( .INP(add_sum[3]), .ZN(n246) );
  NAND4X0 U822 ( .IN1(n446), .IN2(n521), .IN3(n479), .IN4(n522), .QN(n512) );
  OA222X1 U823 ( .IN1(n448), .IN2(n342), .IN3(n424), .IN4(n256), .IN5(n436), 
        .IN6(n259), .Q(n522) );
  OA21X1 U824 ( .IN1(n504), .IN2(n523), .IN3(n479), .Q(n424) );
  INVX0 U825 ( .INP(add_sum[10]), .ZN(n342) );
  OA21X1 U826 ( .IN1(n77), .IN2(n523), .IN3(n436), .Q(n448) );
  OA21X1 U827 ( .IN1(n504), .IN2(n74), .IN3(n479), .Q(n436) );
  NAND2X0 U828 ( .IN1(add_sum[11]), .IN2(n457), .QN(n521) );
  INVX0 U829 ( .INP(n503), .ZN(n457) );
  OA21X1 U830 ( .IN1(n77), .IN2(n74), .IN3(n479), .Q(n503) );
  AND3X1 U831 ( .IN1(n465), .IN2(n328), .IN3(n464), .Q(n446) );
  AND2X1 U832 ( .IN1(n477), .IN2(n330), .Q(n464) );
  AND3X1 U833 ( .IN1(n482), .IN2(n331), .IN3(n480), .Q(n477) );
  AND2X1 U834 ( .IN1(n485), .IN2(n324), .Q(n480) );
  INVX0 U835 ( .INP(add_sum[19]), .ZN(n324) );
  NOR4X0 U836 ( .IN1(n355), .IN2(add_sum[20]), .IN3(add_sum[21]), .IN4(
        add_sum[22]), .QN(n485) );
  AO21X1 U837 ( .IN1(n524), .IN2(n525), .IN3(add_sum[23]), .Q(n355) );
  NOR4X0 U838 ( .IN1(n526), .IN2(n527), .IN3(add_sum[19]), .IN4(add_sum[16]), 
        .QN(n525) );
  NAND3X0 U839 ( .IN1(n321), .IN2(n320), .IN3(n323), .QN(n527) );
  INVX0 U840 ( .INP(add_sum[20]), .ZN(n323) );
  INVX0 U841 ( .INP(add_sum[22]), .ZN(n320) );
  INVX0 U842 ( .INP(add_sum[21]), .ZN(n321) );
  NAND4X0 U843 ( .IN1(n256), .IN2(n259), .IN3(n250), .IN4(n528), .QN(n526) );
  NOR2X0 U844 ( .IN1(add_sum[6]), .IN2(add_sum[3]), .QN(n528) );
  INVX0 U845 ( .INP(add_sum[7]), .ZN(n250) );
  INVX0 U846 ( .INP(add_sum[9]), .ZN(n259) );
  INVX0 U847 ( .INP(add_sum[8]), .ZN(n256) );
  NOR4X0 U848 ( .IN1(n529), .IN2(n530), .IN3(add_sum[10]), .IN4(add_sum[0]), 
        .QN(n524) );
  NAND3X0 U849 ( .IN1(n328), .IN2(n330), .IN3(n358), .QN(n530) );
  INVX0 U850 ( .INP(add_sum[11]), .ZN(n358) );
  INVX0 U851 ( .INP(add_sum[15]), .ZN(n330) );
  NAND4X0 U852 ( .IN1(n361), .IN2(n294), .IN3(n482), .IN4(n465), .QN(n529) );
  NOR2X0 U853 ( .IN1(add_sum[1]), .IN2(add_sum[2]), .QN(n294) );
  NOR2X0 U854 ( .IN1(add_sum[4]), .IN2(add_sum[5]), .QN(n361) );
  INVX0 U855 ( .INP(add_sum[16]), .ZN(n331) );
  INVX0 U856 ( .INP(n505), .ZN(n482) );
  NAND2X0 U857 ( .IN1(n329), .IN2(n325), .QN(n505) );
  INVX0 U858 ( .INP(add_sum[18]), .ZN(n325) );
  INVX0 U859 ( .INP(add_sum[17]), .ZN(n329) );
  INVX0 U860 ( .INP(add_sum[12]), .ZN(n328) );
  NOR2X0 U861 ( .IN1(add_sum[13]), .IN2(add_sum[14]), .QN(n465) );
  OA21X1 U862 ( .IN1(n531), .IN2(n491), .IN3(n366), .Q(add_exception1) );
  XNOR2X1 U863 ( .IN1(add_sign_b), .IN2(add_sign_a), .Q(n366) );
  AND2X1 U864 ( .IN1(n490), .IN2(n67), .Q(n491) );
  AND3X1 U865 ( .IN1(n479), .IN2(n70), .IN3(n487), .Q(n490) );
  NOR2X0 U866 ( .IN1(N841), .IN2(n73), .QN(n487) );
  INVX0 U867 ( .INP(n412), .ZN(n479) );
  NAND2X0 U868 ( .IN1(n517), .IN2(n81), .QN(n412) );
  NOR3X0 U869 ( .IN1(add_new_exponent[6]), .IN2(n87), .IN3(n82), .QN(n517) );
  NOR4X0 U870 ( .IN1(n532), .IN2(n504), .IN3(n81), .IN4(n523), .QN(n531) );
  INVX0 U871 ( .INP(n506), .ZN(n523) );
  NOR2X0 U872 ( .IN1(n67), .IN2(n74), .QN(n506) );
  NAND2X0 U873 ( .IN1(N841), .IN2(n69), .QN(n504) );
  NAND3X0 U874 ( .IN1(n86), .IN2(add_new_exponent[7]), .IN3(n83), .QN(n532) );
endmodule


module booth4_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(SUM[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module booth4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n23), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  NAND2X0 U1 ( .IN1(A[46]), .IN2(carry[46]), .QN(n2) );
  XOR3X1 U2 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X1 U3 ( .IN1(A[46]), .IN2(B[46]), .QN(n1) );
  NAND2X0 U4 ( .IN1(B[46]), .IN2(carry[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[47]) );
  XOR2X1 U6 ( .IN1(A[47]), .IN2(B[47]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[47]), .Q(SUM[47]) );
  NAND2X0 U8 ( .IN1(A[47]), .IN2(B[47]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[47]), .IN2(carry[47]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[47]), .IN2(carry[47]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[48]) );
  XOR3X2 U12 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U13 ( .IN1(A[38]), .IN2(B[38]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[38]), .IN2(carry[38]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[38]), .IN2(carry[38]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[39]) );
  XOR2X1 U17 ( .IN1(A[39]), .IN2(B[39]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U19 ( .IN1(A[39]), .IN2(B[39]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[39]), .IN2(carry[39]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[39]), .IN2(carry[39]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[40]) );
  DELLN2X2 U23 ( .INP(carry[41]), .Z(n15) );
  XOR3X2 U24 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  NAND2X0 U25 ( .IN1(A[40]), .IN2(B[40]), .QN(n16) );
  NAND2X0 U26 ( .IN1(A[40]), .IN2(carry[40]), .QN(n17) );
  NAND2X0 U27 ( .IN1(B[40]), .IN2(carry[40]), .QN(n18) );
  NAND3X0 U28 ( .IN1(n18), .IN2(n17), .IN3(n16), .QN(carry[41]) );
  XOR2X1 U29 ( .IN1(A[41]), .IN2(B[41]), .Q(n19) );
  XOR2X1 U30 ( .IN1(n19), .IN2(n15), .Q(SUM[41]) );
  NAND2X0 U31 ( .IN1(A[41]), .IN2(B[41]), .QN(n20) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(carry[41]), .QN(n21) );
  NAND2X0 U33 ( .IN1(B[41]), .IN2(carry[41]), .QN(n22) );
  NAND3X0 U34 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(carry[42]) );
  AND2X1 U35 ( .IN1(A[26]), .IN2(B[26]), .Q(n23) );
  XOR2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n26), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX2 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX2 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  XOR3X1 U1 ( .IN1(carry[43]), .IN2(B[43]), .IN3(A[43]), .Q(SUM[43]) );
  NAND2X1 U2 ( .IN1(A[43]), .IN2(carry[43]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[43]), .IN2(carry[43]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[43]), .IN2(A[43]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[44]) );
  XOR3X1 U6 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U7 ( .IN1(A[41]), .IN2(B[41]), .IN3(carry[41]), .Q(SUM[41]) );
  NAND2X1 U8 ( .IN1(A[41]), .IN2(B[41]), .QN(n4) );
  NAND2X1 U9 ( .IN1(A[41]), .IN2(carry[41]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[41]), .IN2(carry[41]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[42]) );
  XOR2X1 U12 ( .IN1(A[42]), .IN2(B[42]), .Q(n7) );
  XOR2X1 U13 ( .IN1(n7), .IN2(carry[42]), .Q(SUM[42]) );
  NAND2X0 U14 ( .IN1(A[42]), .IN2(B[42]), .QN(n8) );
  NAND2X0 U15 ( .IN1(A[42]), .IN2(carry[42]), .QN(n9) );
  NAND2X0 U16 ( .IN1(B[42]), .IN2(carry[42]), .QN(n10) );
  NAND3X0 U17 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[43]) );
  DELLN2X2 U18 ( .INP(carry[45]), .Z(n11) );
  XOR3X2 U19 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(B[44]), .QN(n12) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(carry[44]), .QN(n13) );
  NAND2X0 U22 ( .IN1(B[44]), .IN2(carry[44]), .QN(n14) );
  NAND3X0 U23 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[45]) );
  XOR2X1 U24 ( .IN1(A[45]), .IN2(B[45]), .Q(n15) );
  XOR2X1 U25 ( .IN1(n15), .IN2(n11), .Q(SUM[45]) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(B[45]), .QN(n16) );
  NAND2X0 U27 ( .IN1(A[45]), .IN2(carry[45]), .QN(n17) );
  NAND2X0 U28 ( .IN1(B[45]), .IN2(carry[45]), .QN(n18) );
  NAND3X0 U29 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[46]) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U32 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U33 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[48]) );
  XOR2X1 U34 ( .IN1(A[48]), .IN2(B[48]), .Q(n22) );
  XOR2X1 U35 ( .IN1(n22), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(B[48]), .QN(n23) );
  NAND2X0 U37 ( .IN1(A[48]), .IN2(carry[48]), .QN(n24) );
  NAND2X0 U38 ( .IN1(B[48]), .IN2(carry[48]), .QN(n25) );
  NAND3X0 U39 ( .IN1(n23), .IN2(n24), .IN3(n25), .QN(carry[49]) );
  AND2X1 U40 ( .IN1(A[26]), .IN2(B[26]), .Q(n26) );
  XOR2X1 U41 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth4_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[7]), .IN2(A[7]), .Q(SUM[7]) );
endmodule


module booth4 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_sign_a, add_sign_b, 
        add_updated_sum, add_updated_exponent, add_final_exponent_o, 
        add_final_sum_o, add_exception3_o, add_new_sign2, add_new_sign3, 
        add_exception1, add_exception2, add_exception12, add_exception22, s, 
        s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [24:0] add_updated_sum;
  input [7:0] add_updated_exponent;
  output [7:0] add_final_exponent_o;
  output [24:0] add_final_sum_o;
  input clk, reset, new_sign, add_sign_a, add_sign_b, add_new_sign2,
         add_exception1, add_exception2, s;
  output new_sign2, add_exception3_o, add_new_sign3, add_exception12,
         add_exception22, s2;
  wire   N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, add_exception3, N142, N143, N144, N145,
         N146, N147, N148, N149, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n4, n5, n6, n7, n8, n9, n10, n11, n12, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   [24:0] add_final_sum;
  wire   [7:0] add_final_exponent;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[22] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n105), .Q(new_sign2)
         );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n105), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n105), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n105), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n104), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n103), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n102), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n101), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n100), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n99), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n99), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n99), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n40), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n46), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n52), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n58), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n64), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n70), .CLK(clk), .RSTB(n99), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n98), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n98), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n97), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n97), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n97), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n97), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n97), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n6), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n12), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n42), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n48), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n54), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n60), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n66), .CLK(clk), .RSTB(n97), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n72), .CLK(clk), .RSTB(n96), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n96), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n96), 
        .Q(new_exponent2[0]) );
  DFFARX1 add_exception12_reg ( .D(add_exception1), .CLK(clk), .RSTB(n96), .Q(
        add_exception12) );
  DFFARX1 add_exception22_reg ( .D(add_exception2), .CLK(clk), .RSTB(n95), .Q(
        add_exception22) );
  DFFARX1 add_exception3_o_reg ( .D(add_exception3), .CLK(clk), .RSTB(n95), 
        .Q(add_exception3_o) );
  DFFARX1 \add_final_sum_o_reg[24]  ( .D(add_final_sum[24]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[24]) );
  DFFARX1 \add_final_sum_o_reg[23]  ( .D(add_final_sum[23]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[23]) );
  DFFARX1 \add_final_sum_o_reg[22]  ( .D(add_final_sum[22]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[22]) );
  DFFARX1 \add_final_sum_o_reg[21]  ( .D(add_final_sum[21]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[21]) );
  DFFARX1 \add_final_sum_o_reg[20]  ( .D(add_final_sum[20]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[20]) );
  DFFARX1 \add_final_sum_o_reg[19]  ( .D(add_final_sum[19]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[19]) );
  DFFARX1 \add_final_sum_o_reg[18]  ( .D(add_final_sum[18]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[18]) );
  DFFARX1 \add_final_sum_o_reg[17]  ( .D(add_final_sum[17]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[17]) );
  DFFARX1 \add_final_sum_o_reg[16]  ( .D(add_final_sum[16]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[16]) );
  DFFARX1 \add_final_sum_o_reg[15]  ( .D(add_final_sum[15]), .CLK(clk), .RSTB(
        n95), .Q(add_final_sum_o[15]) );
  DFFARX1 \add_final_sum_o_reg[14]  ( .D(add_final_sum[14]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[14]) );
  DFFARX1 \add_final_sum_o_reg[13]  ( .D(add_final_sum[13]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[13]) );
  DFFARX1 \add_final_sum_o_reg[12]  ( .D(add_final_sum[12]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[12]) );
  DFFARX1 \add_final_sum_o_reg[11]  ( .D(add_final_sum[11]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[11]) );
  DFFARX1 \add_final_sum_o_reg[10]  ( .D(add_final_sum[10]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[10]) );
  DFFARX1 \add_final_sum_o_reg[9]  ( .D(add_final_sum[9]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[9]) );
  DFFARX1 \add_final_sum_o_reg[8]  ( .D(add_final_sum[8]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[8]) );
  DFFARX1 \add_final_sum_o_reg[7]  ( .D(add_final_sum[7]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[7]) );
  DFFARX1 \add_final_sum_o_reg[6]  ( .D(add_final_sum[6]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[6]) );
  DFFARX1 \add_final_sum_o_reg[5]  ( .D(add_final_sum[5]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[5]) );
  DFFARX1 \add_final_sum_o_reg[4]  ( .D(add_final_sum[4]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[4]) );
  DFFARX1 \add_final_sum_o_reg[3]  ( .D(add_final_sum[3]), .CLK(clk), .RSTB(
        n94), .Q(add_final_sum_o[3]) );
  DFFARX1 \add_final_sum_o_reg[2]  ( .D(add_final_sum[2]), .CLK(clk), .RSTB(
        n93), .Q(add_final_sum_o[2]) );
  DFFARX1 \add_final_sum_o_reg[1]  ( .D(add_final_sum[1]), .CLK(clk), .RSTB(
        n93), .Q(add_final_sum_o[1]) );
  DFFARX1 \add_final_sum_o_reg[0]  ( .D(add_final_sum[0]), .CLK(clk), .RSTB(
        n93), .Q(add_final_sum_o[0]) );
  DFFARX1 \add_final_exponent_o_reg[7]  ( .D(add_final_exponent[7]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[7]) );
  DFFARX1 \add_final_exponent_o_reg[6]  ( .D(add_final_exponent[6]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[6]) );
  DFFARX1 \add_final_exponent_o_reg[5]  ( .D(add_final_exponent[5]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[5]) );
  DFFARX1 \add_final_exponent_o_reg[4]  ( .D(add_final_exponent[4]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[4]) );
  DFFARX1 \add_final_exponent_o_reg[3]  ( .D(add_final_exponent[3]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[3]) );
  DFFARX1 \add_final_exponent_o_reg[2]  ( .D(add_final_exponent[2]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[2]) );
  DFFARX1 \add_final_exponent_o_reg[1]  ( .D(add_final_exponent[1]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[1]) );
  DFFARX1 \add_final_exponent_o_reg[0]  ( .D(add_final_exponent[0]), .CLK(clk), 
        .RSTB(n93), .Q(add_final_exponent_o[0]) );
  DFFARX1 add_new_sign3_reg ( .D(add_new_sign2), .CLK(clk), .RSTB(n93), .Q(
        add_new_sign3) );
  AO222X1 U17 ( .IN1(N31), .IN2(n89), .IN3(N82), .IN4(n86), .IN5(
        product_shift[9]), .IN6(n84), .Q(product2[9]) );
  AO222X1 U18 ( .IN1(N30), .IN2(n89), .IN3(N81), .IN4(n86), .IN5(
        product_shift[8]), .IN6(n15), .Q(product2[8]) );
  AO222X1 U19 ( .IN1(N29), .IN2(n89), .IN3(N80), .IN4(n86), .IN5(
        product_shift[7]), .IN6(n15), .Q(product2[7]) );
  AO222X1 U20 ( .IN1(N28), .IN2(n89), .IN3(N79), .IN4(n86), .IN5(
        product_shift[6]), .IN6(n15), .Q(product2[6]) );
  AO222X1 U21 ( .IN1(N27), .IN2(n89), .IN3(N78), .IN4(n86), .IN5(
        product_shift[5]), .IN6(n15), .Q(product2[5]) );
  AO222X1 U22 ( .IN1(N72), .IN2(n89), .IN3(N123), .IN4(n86), .IN5(
        product_shift[49]), .IN6(n15), .Q(product2[50]) );
  AO222X1 U23 ( .IN1(N26), .IN2(n89), .IN3(N77), .IN4(n86), .IN5(
        product_shift[4]), .IN6(n84), .Q(product2[4]) );
  AO222X1 U24 ( .IN1(N71), .IN2(n89), .IN3(N122), .IN4(n86), .IN5(
        product_shift[49]), .IN6(n85), .Q(product2[49]) );
  AO222X1 U25 ( .IN1(N70), .IN2(n89), .IN3(N121), .IN4(n86), .IN5(
        product_shift[48]), .IN6(n15), .Q(product2[48]) );
  AO222X1 U26 ( .IN1(N69), .IN2(n89), .IN3(N120), .IN4(n86), .IN5(
        product_shift[47]), .IN6(n85), .Q(product2[47]) );
  AO222X1 U27 ( .IN1(N68), .IN2(n89), .IN3(N119), .IN4(n86), .IN5(
        product_shift[46]), .IN6(n15), .Q(product2[46]) );
  AO222X1 U28 ( .IN1(N67), .IN2(n89), .IN3(N118), .IN4(n86), .IN5(
        product_shift[45]), .IN6(n15), .Q(product2[45]) );
  AO222X1 U29 ( .IN1(N66), .IN2(n90), .IN3(N117), .IN4(n87), .IN5(
        product_shift[44]), .IN6(n85), .Q(product2[44]) );
  AO222X1 U30 ( .IN1(N65), .IN2(n90), .IN3(N116), .IN4(n87), .IN5(
        product_shift[43]), .IN6(n85), .Q(product2[43]) );
  AO222X1 U31 ( .IN1(N64), .IN2(n90), .IN3(N115), .IN4(n87), .IN5(
        product_shift[42]), .IN6(n85), .Q(product2[42]) );
  AO222X1 U32 ( .IN1(N63), .IN2(n90), .IN3(N114), .IN4(n87), .IN5(
        product_shift[41]), .IN6(n85), .Q(product2[41]) );
  AO222X1 U33 ( .IN1(N62), .IN2(n90), .IN3(N113), .IN4(n87), .IN5(
        product_shift[40]), .IN6(n85), .Q(product2[40]) );
  AO222X1 U34 ( .IN1(N25), .IN2(n90), .IN3(N76), .IN4(n87), .IN5(
        product_shift[3]), .IN6(n85), .Q(product2[3]) );
  AO222X1 U35 ( .IN1(N61), .IN2(n90), .IN3(N112), .IN4(n87), .IN5(
        product_shift[39]), .IN6(n85), .Q(product2[39]) );
  AO222X1 U36 ( .IN1(N60), .IN2(n90), .IN3(N111), .IN4(n87), .IN5(
        product_shift[38]), .IN6(n85), .Q(product2[38]) );
  AO222X1 U37 ( .IN1(N59), .IN2(n90), .IN3(N110), .IN4(n87), .IN5(
        product_shift[37]), .IN6(n85), .Q(product2[37]) );
  AO222X1 U38 ( .IN1(N58), .IN2(n90), .IN3(N109), .IN4(n87), .IN5(
        product_shift[36]), .IN6(n85), .Q(product2[36]) );
  AO222X1 U39 ( .IN1(N57), .IN2(n90), .IN3(N108), .IN4(n87), .IN5(n4), .IN6(
        n85), .Q(product2[35]) );
  AO222X1 U40 ( .IN1(N56), .IN2(n90), .IN3(N107), .IN4(n87), .IN5(n8), .IN6(
        n85), .Q(product2[34]) );
  AO222X1 U41 ( .IN1(N55), .IN2(n91), .IN3(N106), .IN4(n88), .IN5(n38), .IN6(
        n85), .Q(product2[33]) );
  AO222X1 U42 ( .IN1(N54), .IN2(n91), .IN3(N105), .IN4(n88), .IN5(n44), .IN6(
        n15), .Q(product2[32]) );
  AO222X1 U43 ( .IN1(N53), .IN2(n91), .IN3(N104), .IN4(n88), .IN5(n50), .IN6(
        n15), .Q(product2[31]) );
  AO222X1 U44 ( .IN1(N52), .IN2(n91), .IN3(N103), .IN4(n88), .IN5(n56), .IN6(
        n15), .Q(product2[30]) );
  AO222X1 U45 ( .IN1(N24), .IN2(n91), .IN3(N75), .IN4(n88), .IN5(
        product_shift[2]), .IN6(n15), .Q(product2[2]) );
  AO222X1 U46 ( .IN1(N51), .IN2(n91), .IN3(N102), .IN4(n88), .IN5(n62), .IN6(
        n15), .Q(product2[29]) );
  AO222X1 U47 ( .IN1(N50), .IN2(n91), .IN3(N101), .IN4(n88), .IN5(n68), .IN6(
        n15), .Q(product2[28]) );
  AO222X1 U48 ( .IN1(N49), .IN2(n91), .IN3(N100), .IN4(n88), .IN5(n74), .IN6(
        n15), .Q(product2[27]) );
  AO222X1 U49 ( .IN1(N48), .IN2(n91), .IN3(N99), .IN4(n88), .IN5(n76), .IN6(
        n15), .Q(product2[26]) );
  AO222X1 U50 ( .IN1(N47), .IN2(n91), .IN3(N98), .IN4(n88), .IN5(
        product_shift[25]), .IN6(n15), .Q(product2[25]) );
  AO222X1 U51 ( .IN1(N46), .IN2(n91), .IN3(N97), .IN4(n88), .IN5(
        product_shift[24]), .IN6(n15), .Q(product2[24]) );
  AO222X1 U52 ( .IN1(N45), .IN2(n91), .IN3(N96), .IN4(n88), .IN5(
        product_shift[23]), .IN6(n84), .Q(product2[23]) );
  AO222X1 U54 ( .IN1(N43), .IN2(n92), .IN3(N94), .IN4(n14), .IN5(
        product_shift[21]), .IN6(n84), .Q(product2[21]) );
  AO222X1 U55 ( .IN1(N42), .IN2(n92), .IN3(N93), .IN4(n14), .IN5(
        product_shift[20]), .IN6(n84), .Q(product2[20]) );
  AO222X1 U56 ( .IN1(N23), .IN2(n92), .IN3(N74), .IN4(n88), .IN5(n84), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U57 ( .IN1(N41), .IN2(n92), .IN3(N92), .IN4(n14), .IN5(
        product_shift[19]), .IN6(n84), .Q(product2[19]) );
  AO222X1 U58 ( .IN1(N40), .IN2(n92), .IN3(N91), .IN4(n14), .IN5(
        product_shift[18]), .IN6(n84), .Q(product2[18]) );
  AO222X1 U59 ( .IN1(N39), .IN2(n92), .IN3(N90), .IN4(n14), .IN5(
        product_shift[17]), .IN6(n84), .Q(product2[17]) );
  AO222X1 U60 ( .IN1(N38), .IN2(n92), .IN3(N89), .IN4(n14), .IN5(
        product_shift[16]), .IN6(n84), .Q(product2[16]) );
  AO222X1 U61 ( .IN1(N37), .IN2(n92), .IN3(N88), .IN4(n14), .IN5(
        product_shift[15]), .IN6(n84), .Q(product2[15]) );
  AO222X1 U62 ( .IN1(N36), .IN2(n92), .IN3(N87), .IN4(n14), .IN5(
        product_shift[14]), .IN6(n84), .Q(product2[14]) );
  AO222X1 U63 ( .IN1(N35), .IN2(n92), .IN3(N86), .IN4(n14), .IN5(
        product_shift[13]), .IN6(n84), .Q(product2[13]) );
  AO222X1 U64 ( .IN1(N34), .IN2(n92), .IN3(N85), .IN4(n14), .IN5(
        product_shift[12]), .IN6(n84), .Q(product2[12]) );
  AO222X1 U65 ( .IN1(N33), .IN2(n92), .IN3(N84), .IN4(n86), .IN5(
        product_shift[11]), .IN6(n84), .Q(product2[11]) );
  AO222X1 U66 ( .IN1(N32), .IN2(n92), .IN3(N83), .IN4(n87), .IN5(
        product_shift[10]), .IN6(n85), .Q(product2[10]) );
  XOR2X1 U68 ( .IN1(n106), .IN2(product_shift[1]), .Q(n15) );
  AND2X1 U69 ( .IN1(product_shift[1]), .IN2(n106), .Q(n14) );
  AO222X1 U70 ( .IN1(N160), .IN2(n78), .IN3(add_updated_sum[10]), .IN4(n80), 
        .IN5(add_updated_sum[9]), .IN6(n81), .Q(add_final_sum[9]) );
  AO222X1 U71 ( .IN1(N159), .IN2(n78), .IN3(add_updated_sum[9]), .IN4(n80), 
        .IN5(add_updated_sum[8]), .IN6(n81), .Q(add_final_sum[8]) );
  AO222X1 U72 ( .IN1(N158), .IN2(n78), .IN3(add_updated_sum[8]), .IN4(n80), 
        .IN5(add_updated_sum[7]), .IN6(n81), .Q(add_final_sum[7]) );
  AO222X1 U73 ( .IN1(N157), .IN2(n78), .IN3(add_updated_sum[7]), .IN4(n80), 
        .IN5(add_updated_sum[6]), .IN6(n81), .Q(add_final_sum[6]) );
  AO222X1 U74 ( .IN1(N156), .IN2(n78), .IN3(add_updated_sum[6]), .IN4(n80), 
        .IN5(add_updated_sum[5]), .IN6(n81), .Q(add_final_sum[5]) );
  AO222X1 U75 ( .IN1(N155), .IN2(n78), .IN3(add_updated_sum[5]), .IN4(n80), 
        .IN5(add_updated_sum[4]), .IN6(n81), .Q(add_final_sum[4]) );
  AO222X1 U76 ( .IN1(N154), .IN2(n78), .IN3(add_updated_sum[4]), .IN4(n80), 
        .IN5(add_updated_sum[3]), .IN6(n81), .Q(add_final_sum[3]) );
  AO222X1 U77 ( .IN1(N153), .IN2(n78), .IN3(add_updated_sum[3]), .IN4(n80), 
        .IN5(add_updated_sum[2]), .IN6(n81), .Q(add_final_sum[2]) );
  AO22X1 U78 ( .IN1(add_updated_sum[24]), .IN2(n107), .IN3(N175), .IN4(n78), 
        .Q(add_final_sum[24]) );
  AO222X1 U79 ( .IN1(N174), .IN2(n78), .IN3(add_updated_sum[24]), .IN4(n80), 
        .IN5(add_updated_sum[23]), .IN6(n81), .Q(add_final_sum[23]) );
  AO222X1 U80 ( .IN1(N173), .IN2(n78), .IN3(n80), .IN4(add_updated_sum[23]), 
        .IN5(add_updated_sum[22]), .IN6(n81), .Q(add_final_sum[22]) );
  AO222X1 U81 ( .IN1(N172), .IN2(n78), .IN3(add_updated_sum[22]), .IN4(n80), 
        .IN5(add_updated_sum[21]), .IN6(n81), .Q(add_final_sum[21]) );
  AO222X1 U82 ( .IN1(N171), .IN2(n79), .IN3(add_updated_sum[21]), .IN4(n80), 
        .IN5(add_updated_sum[20]), .IN6(n81), .Q(add_final_sum[20]) );
  AO222X1 U83 ( .IN1(N152), .IN2(n79), .IN3(add_updated_sum[2]), .IN4(n109), 
        .IN5(add_updated_sum[1]), .IN6(n82), .Q(add_final_sum[1]) );
  AO222X1 U84 ( .IN1(N170), .IN2(n79), .IN3(add_updated_sum[20]), .IN4(n109), 
        .IN5(add_updated_sum[19]), .IN6(n82), .Q(add_final_sum[19]) );
  AO222X1 U85 ( .IN1(N169), .IN2(n79), .IN3(add_updated_sum[19]), .IN4(n109), 
        .IN5(add_updated_sum[18]), .IN6(n82), .Q(add_final_sum[18]) );
  AO222X1 U86 ( .IN1(N168), .IN2(n79), .IN3(add_updated_sum[18]), .IN4(n109), 
        .IN5(add_updated_sum[17]), .IN6(n82), .Q(add_final_sum[17]) );
  AO222X1 U87 ( .IN1(N167), .IN2(n79), .IN3(add_updated_sum[17]), .IN4(n109), 
        .IN5(add_updated_sum[16]), .IN6(n82), .Q(add_final_sum[16]) );
  AO222X1 U88 ( .IN1(N166), .IN2(n79), .IN3(add_updated_sum[16]), .IN4(n109), 
        .IN5(add_updated_sum[15]), .IN6(n82), .Q(add_final_sum[15]) );
  AO222X1 U89 ( .IN1(N165), .IN2(n79), .IN3(add_updated_sum[15]), .IN4(n109), 
        .IN5(add_updated_sum[14]), .IN6(n82), .Q(add_final_sum[14]) );
  AO222X1 U90 ( .IN1(N164), .IN2(n79), .IN3(add_updated_sum[14]), .IN4(n109), 
        .IN5(add_updated_sum[13]), .IN6(n82), .Q(add_final_sum[13]) );
  AO222X1 U91 ( .IN1(N163), .IN2(n79), .IN3(add_updated_sum[13]), .IN4(n109), 
        .IN5(add_updated_sum[12]), .IN6(n82), .Q(add_final_sum[12]) );
  AO222X1 U92 ( .IN1(N162), .IN2(n79), .IN3(add_updated_sum[12]), .IN4(n80), 
        .IN5(add_updated_sum[11]), .IN6(n82), .Q(add_final_sum[11]) );
  AO222X1 U93 ( .IN1(N161), .IN2(n79), .IN3(add_updated_sum[11]), .IN4(n80), 
        .IN5(add_updated_sum[10]), .IN6(n82), .Q(add_final_sum[10]) );
  AO222X1 U94 ( .IN1(N151), .IN2(n78), .IN3(add_updated_sum[1]), .IN4(n80), 
        .IN5(add_updated_sum[0]), .IN6(n82), .Q(add_final_sum[0]) );
  AO22X1 U95 ( .IN1(add_updated_exponent[7]), .IN2(n83), .IN3(N149), .IN4(n19), 
        .Q(add_final_exponent[7]) );
  AO22X1 U96 ( .IN1(add_updated_exponent[6]), .IN2(n83), .IN3(N148), .IN4(n19), 
        .Q(add_final_exponent[6]) );
  AO22X1 U97 ( .IN1(add_updated_exponent[5]), .IN2(n83), .IN3(N147), .IN4(n19), 
        .Q(add_final_exponent[5]) );
  AO22X1 U98 ( .IN1(add_updated_exponent[4]), .IN2(n83), .IN3(N146), .IN4(n19), 
        .Q(add_final_exponent[4]) );
  AO22X1 U99 ( .IN1(add_updated_exponent[3]), .IN2(n83), .IN3(N145), .IN4(n19), 
        .Q(add_final_exponent[3]) );
  AO22X1 U100 ( .IN1(add_updated_exponent[2]), .IN2(n83), .IN3(N144), .IN4(n19), .Q(add_final_exponent[2]) );
  AO22X1 U101 ( .IN1(add_updated_exponent[1]), .IN2(n83), .IN3(N143), .IN4(n19), .Q(add_final_exponent[1]) );
  AO22X1 U102 ( .IN1(add_updated_exponent[0]), .IN2(n83), .IN3(N142), .IN4(n19), .Q(add_final_exponent[0]) );
  NAND3X0 U103 ( .IN1(n20), .IN2(n111), .IN3(n21), .QN(n17) );
  NAND3X0 U104 ( .IN1(n21), .IN2(n20), .IN3(add_updated_sum[0]), .QN(n18) );
  XNOR2X1 U105 ( .IN1(add_sign_b), .IN2(add_sign_a), .Q(n21) );
  OA22X1 U106 ( .IN1(n23), .IN2(n24), .IN3(n25), .IN4(n26), .Q(n22) );
  NAND4X0 U107 ( .IN1(add_updated_exponent[0]), .IN2(add_updated_exponent[1]), 
        .IN3(add_updated_exponent[2]), .IN4(add_updated_exponent[3]), .QN(n26)
         );
  NAND4X0 U108 ( .IN1(add_updated_exponent[4]), .IN2(add_updated_exponent[5]), 
        .IN3(add_updated_exponent[6]), .IN4(add_updated_exponent[7]), .QN(n25)
         );
  OR4X1 U109 ( .IN1(n27), .IN2(add_updated_exponent[0]), .IN3(
        add_updated_exponent[1]), .IN4(add_updated_exponent[2]), .Q(n24) );
  AND4X1 U110 ( .IN1(n28), .IN2(n29), .IN3(n30), .IN4(n31), .Q(n27) );
  NOR4X0 U111 ( .IN1(n32), .IN2(add_updated_sum[4]), .IN3(add_updated_sum[6]), 
        .IN4(add_updated_sum[5]), .QN(n31) );
  OR3X1 U112 ( .IN1(add_updated_sum[8]), .IN2(add_updated_sum[9]), .IN3(
        add_updated_sum[7]), .Q(n32) );
  NOR4X0 U113 ( .IN1(n33), .IN2(add_updated_sum[1]), .IN3(add_updated_sum[21]), 
        .IN4(add_updated_sum[20]), .QN(n30) );
  OR3X1 U114 ( .IN1(add_updated_sum[2]), .IN2(add_updated_sum[3]), .IN3(
        add_updated_sum[22]), .Q(n33) );
  NOR4X0 U115 ( .IN1(n34), .IN2(add_updated_sum[14]), .IN3(add_updated_sum[16]), .IN4(add_updated_sum[15]), .QN(n29) );
  OR3X1 U116 ( .IN1(add_updated_sum[18]), .IN2(add_updated_sum[19]), .IN3(
        add_updated_sum[17]), .Q(n34) );
  NOR4X0 U117 ( .IN1(n35), .IN2(add_updated_sum[11]), .IN3(add_updated_sum[13]), .IN4(add_updated_sum[12]), .QN(n28) );
  OR2X1 U118 ( .IN1(add_updated_sum[0]), .IN2(add_updated_sum[10]), .Q(n35) );
  OR4X1 U119 ( .IN1(add_updated_exponent[3]), .IN2(add_updated_exponent[4]), 
        .IN3(n36), .IN4(add_updated_exponent[5]), .Q(n23) );
  OR2X1 U120 ( .IN1(add_updated_exponent[7]), .IN2(add_updated_exponent[6]), 
        .Q(n36) );
  booth4_DW01_inc_0 add_194 ( .A({1'b0, add_updated_sum[24:1]}), .SUM({N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151}) );
  booth4_DW01_add_0 add_98 ( .A({product_shift[49], product_shift[49:36], n4, 
        n8, n38, n44, n50, n56, n62, n68, n74, n76, product_shift[25:0]}), .B(
        {combined_negative_b[24:9], n6, n12, n42, n48, n54, n60, n66, n72, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N123, N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96, SYNOPSYS_UNCONNECTED__0, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth4_DW01_add_1 add_91 ( .A({product_shift[49], product_shift[49:35], n8, 
        n38, n44, n50, n56, n62, n68, n74, n76, product_shift[25:0]}), .B({
        combined_b[24:8], n10, n40, n46, n52, n58, n64, n70, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, SYNOPSYS_UNCONNECTED__2, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, SYNOPSYS_UNCONNECTED__3}) );
  booth4_DW01_inc_1 r69 ( .A(add_updated_exponent), .SUM({N149, N148, N147, 
        N146, N145, N144, N143, N142}) );
  NBUFFX2 U3 ( .INP(product_shift[35]), .Z(n4) );
  INVX0 U4 ( .INP(combined_negative_b[8]), .ZN(n5) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  INVX0 U6 ( .INP(product_shift[34]), .ZN(n7) );
  INVX0 U7 ( .INP(n7), .ZN(n8) );
  INVX0 U11 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U12 ( .INP(n9), .ZN(n10) );
  INVX0 U13 ( .INP(combined_negative_b[7]), .ZN(n11) );
  INVX0 U14 ( .INP(n11), .ZN(n12) );
  INVX0 U15 ( .INP(product_shift[33]), .ZN(n37) );
  INVX0 U16 ( .INP(n37), .ZN(n38) );
  INVX0 U53 ( .INP(combined_b[6]), .ZN(n39) );
  INVX0 U67 ( .INP(n39), .ZN(n40) );
  INVX0 U121 ( .INP(combined_negative_b[6]), .ZN(n41) );
  INVX0 U122 ( .INP(n41), .ZN(n42) );
  INVX0 U123 ( .INP(product_shift[32]), .ZN(n43) );
  INVX0 U124 ( .INP(n43), .ZN(n44) );
  INVX0 U125 ( .INP(combined_b[5]), .ZN(n45) );
  INVX0 U126 ( .INP(n45), .ZN(n46) );
  INVX0 U127 ( .INP(combined_negative_b[5]), .ZN(n47) );
  INVX0 U128 ( .INP(n47), .ZN(n48) );
  INVX0 U129 ( .INP(product_shift[31]), .ZN(n49) );
  INVX0 U130 ( .INP(n49), .ZN(n50) );
  INVX0 U131 ( .INP(combined_b[4]), .ZN(n51) );
  INVX0 U132 ( .INP(n51), .ZN(n52) );
  INVX0 U133 ( .INP(combined_negative_b[4]), .ZN(n53) );
  INVX0 U134 ( .INP(n53), .ZN(n54) );
  INVX0 U135 ( .INP(product_shift[30]), .ZN(n55) );
  INVX0 U136 ( .INP(n55), .ZN(n56) );
  INVX0 U137 ( .INP(combined_b[3]), .ZN(n57) );
  INVX0 U138 ( .INP(n57), .ZN(n58) );
  INVX0 U139 ( .INP(combined_negative_b[3]), .ZN(n59) );
  INVX0 U140 ( .INP(n59), .ZN(n60) );
  INVX0 U141 ( .INP(product_shift[29]), .ZN(n61) );
  INVX0 U142 ( .INP(n61), .ZN(n62) );
  INVX0 U143 ( .INP(combined_b[2]), .ZN(n63) );
  INVX0 U144 ( .INP(n63), .ZN(n64) );
  INVX0 U145 ( .INP(combined_negative_b[2]), .ZN(n65) );
  INVX0 U146 ( .INP(n65), .ZN(n66) );
  INVX0 U147 ( .INP(product_shift[28]), .ZN(n67) );
  INVX0 U148 ( .INP(n67), .ZN(n68) );
  INVX0 U149 ( .INP(combined_b[1]), .ZN(n69) );
  INVX0 U150 ( .INP(n69), .ZN(n70) );
  INVX0 U151 ( .INP(combined_negative_b[1]), .ZN(n71) );
  INVX0 U152 ( .INP(n71), .ZN(n72) );
  INVX0 U153 ( .INP(product_shift[27]), .ZN(n73) );
  INVX0 U154 ( .INP(n73), .ZN(n74) );
  NBUFFX2 U155 ( .INP(n109), .Z(n80) );
  NBUFFX2 U156 ( .INP(n16), .Z(n82) );
  NBUFFX2 U157 ( .INP(n16), .Z(n81) );
  NBUFFX2 U158 ( .INP(n108), .Z(n78) );
  NBUFFX2 U159 ( .INP(n108), .Z(n79) );
  NBUFFX2 U160 ( .INP(n16), .Z(n83) );
  NBUFFX2 U161 ( .INP(n77), .Z(n93) );
  NBUFFX2 U162 ( .INP(n77), .Z(n94) );
  NBUFFX2 U163 ( .INP(n77), .Z(n95) );
  NBUFFX2 U164 ( .INP(n77), .Z(n96) );
  NBUFFX2 U165 ( .INP(n77), .Z(n97) );
  NBUFFX2 U166 ( .INP(n77), .Z(n98) );
  NBUFFX2 U167 ( .INP(n77), .Z(n99) );
  NBUFFX2 U168 ( .INP(n77), .Z(n100) );
  NBUFFX2 U169 ( .INP(n77), .Z(n101) );
  NBUFFX2 U170 ( .INP(n77), .Z(n103) );
  NBUFFX2 U171 ( .INP(n77), .Z(n104) );
  NBUFFX2 U172 ( .INP(n77), .Z(n102) );
  NBUFFX2 U173 ( .INP(n77), .Z(n105) );
  NBUFFX2 U174 ( .INP(n13), .Z(n91) );
  NBUFFX2 U175 ( .INP(n13), .Z(n90) );
  NBUFFX2 U176 ( .INP(n13), .Z(n89) );
  NBUFFX2 U177 ( .INP(n13), .Z(n92) );
  NBUFFX2 U178 ( .INP(n15), .Z(n84) );
  NBUFFX2 U179 ( .INP(n15), .Z(n85) );
  NAND2X1 U180 ( .IN1(n18), .IN2(n17), .QN(n19) );
  INVX0 U181 ( .INP(n18), .ZN(n108) );
  INVX0 U182 ( .INP(n17), .ZN(n109) );
  NAND2X1 U183 ( .IN1(n21), .IN2(n20), .QN(n16) );
  NBUFFX2 U184 ( .INP(n14), .Z(n88) );
  NBUFFX2 U185 ( .INP(n14), .Z(n87) );
  NBUFFX2 U186 ( .INP(n14), .Z(n86) );
  INVX0 U187 ( .INP(n21), .ZN(n107) );
  NBUFFX2 U188 ( .INP(reset), .Z(n77) );
  NOR2X0 U189 ( .IN1(n106), .IN2(product_shift[1]), .QN(n13) );
  INVX0 U190 ( .INP(add_updated_sum[0]), .ZN(n111) );
  NAND2X1 U191 ( .IN1(add_updated_sum[23]), .IN2(n110), .QN(n20) );
  INVX0 U192 ( .INP(add_updated_sum[24]), .ZN(n110) );
  NOR2X0 U193 ( .IN1(n22), .IN2(n107), .QN(add_exception3) );
  INVX0 U194 ( .INP(product_shift[0]), .ZN(n106) );
  INVX0 U196 ( .INP(product_shift[26]), .ZN(n75) );
  INVX0 U197 ( .INP(n75), .ZN(n76) );
endmodule


module booth5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n35), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  DELLN2X2 U1 ( .INP(carry[46]), .Z(n1) );
  DELLN1X2 U2 ( .INP(carry[47]), .Z(n12) );
  XOR3X1 U3 ( .IN1(carry[48]), .IN2(B[48]), .IN3(A[48]), .Q(SUM[48]) );
  NAND2X1 U4 ( .IN1(A[48]), .IN2(carry[48]), .QN(n2) );
  NAND2X0 U5 ( .IN1(B[48]), .IN2(carry[48]), .QN(n3) );
  NAND2X1 U6 ( .IN1(B[48]), .IN2(A[48]), .QN(n4) );
  NAND3X0 U7 ( .IN1(n2), .IN2(n4), .IN3(n3), .QN(carry[49]) );
  XOR3X1 U8 ( .IN1(carry[45]), .IN2(B[45]), .IN3(A[45]), .Q(SUM[45]) );
  NAND2X0 U9 ( .IN1(A[45]), .IN2(carry[45]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[45]), .IN2(carry[45]), .QN(n6) );
  NAND2X0 U11 ( .IN1(B[45]), .IN2(A[45]), .QN(n7) );
  NAND3X0 U12 ( .IN1(n5), .IN2(n7), .IN3(n6), .QN(carry[46]) );
  XOR3X1 U13 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U14 ( .IN1(A[42]), .IN2(carry[42]), .QN(n8) );
  NAND2X0 U15 ( .IN1(B[42]), .IN2(carry[42]), .QN(n9) );
  NAND2X0 U16 ( .IN1(B[42]), .IN2(A[42]), .QN(n10) );
  NAND3X0 U17 ( .IN1(n8), .IN2(n10), .IN3(n9), .QN(carry[43]) );
  DELLN2X2 U18 ( .INP(carry[44]), .Z(n11) );
  DELLN2X2 U19 ( .INP(carry[41]), .Z(n13) );
  XOR3X2 U20 ( .IN1(A[46]), .IN2(B[46]), .IN3(n1), .Q(SUM[46]) );
  XOR3X2 U21 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U22 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U23 ( .IN1(A[40]), .IN2(B[40]), .QN(n14) );
  NAND2X0 U24 ( .IN1(A[40]), .IN2(carry[40]), .QN(n15) );
  NAND2X0 U25 ( .IN1(B[40]), .IN2(carry[40]), .QN(n16) );
  NAND3X0 U26 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[41]) );
  XOR2X1 U27 ( .IN1(A[41]), .IN2(B[41]), .Q(n17) );
  XOR2X1 U28 ( .IN1(n17), .IN2(n13), .Q(SUM[41]) );
  NAND2X0 U29 ( .IN1(A[41]), .IN2(B[41]), .QN(n18) );
  NAND2X0 U30 ( .IN1(A[41]), .IN2(carry[41]), .QN(n19) );
  NAND2X0 U31 ( .IN1(B[41]), .IN2(carry[41]), .QN(n20) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[42]) );
  NAND2X0 U33 ( .IN1(A[43]), .IN2(B[43]), .QN(n21) );
  NAND2X0 U34 ( .IN1(A[43]), .IN2(carry[43]), .QN(n22) );
  NAND2X0 U35 ( .IN1(B[43]), .IN2(carry[43]), .QN(n23) );
  NAND3X0 U36 ( .IN1(n22), .IN2(n23), .IN3(n21), .QN(carry[44]) );
  XOR2X1 U37 ( .IN1(A[44]), .IN2(B[44]), .Q(n24) );
  XOR2X1 U38 ( .IN1(n24), .IN2(n11), .Q(SUM[44]) );
  NAND2X0 U39 ( .IN1(A[44]), .IN2(B[44]), .QN(n25) );
  NAND2X0 U40 ( .IN1(A[44]), .IN2(carry[44]), .QN(n26) );
  NAND2X0 U41 ( .IN1(B[44]), .IN2(carry[44]), .QN(n27) );
  NAND3X0 U42 ( .IN1(n26), .IN2(n27), .IN3(n25), .QN(carry[45]) );
  NAND2X0 U43 ( .IN1(A[46]), .IN2(B[46]), .QN(n28) );
  NAND2X0 U44 ( .IN1(A[46]), .IN2(carry[46]), .QN(n29) );
  NAND2X0 U45 ( .IN1(B[46]), .IN2(carry[46]), .QN(n30) );
  NAND3X0 U46 ( .IN1(n28), .IN2(n29), .IN3(n30), .QN(carry[47]) );
  XOR2X1 U47 ( .IN1(A[47]), .IN2(B[47]), .Q(n31) );
  XOR2X1 U48 ( .IN1(n31), .IN2(n12), .Q(SUM[47]) );
  NAND2X0 U49 ( .IN1(A[47]), .IN2(B[47]), .QN(n32) );
  NAND2X0 U50 ( .IN1(A[47]), .IN2(carry[47]), .QN(n33) );
  NAND2X0 U51 ( .IN1(B[47]), .IN2(carry[47]), .QN(n34) );
  NAND3X0 U52 ( .IN1(n33), .IN2(n34), .IN3(n32), .QN(carry[48]) );
  AND2X1 U53 ( .IN1(A[26]), .IN2(B[26]), .Q(n35) );
  XOR2X1 U54 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n24), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X1 U1 ( .IN1(carry[39]), .IN2(B[39]), .IN3(A[39]), .Q(SUM[39]) );
  NAND2X0 U2 ( .IN1(A[39]), .IN2(carry[39]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[39]), .IN2(carry[39]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[39]), .IN2(A[39]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[40]) );
  XOR3X1 U6 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U7 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[50]) );
  DELLN2X2 U11 ( .INP(carry[45]), .Z(n7) );
  INVX0 U12 ( .INP(A[34]), .ZN(n8) );
  INVX0 U13 ( .INP(n8), .ZN(n9) );
  XOR3X1 U14 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U16 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U17 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U18 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U19 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U20 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U21 ( .IN1(n13), .IN2(n7), .Q(SUM[45]) );
  NAND2X0 U22 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U23 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U24 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U25 ( .IN1(n16), .IN2(n15), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U26 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U27 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U28 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U29 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U30 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U31 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U32 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U34 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U35 ( .IN1(n23), .IN2(n22), .IN3(n21), .QN(carry[49]) );
  AND2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(n24) );
  XOR2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth5 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_final_exponent, add_final_sum, 
        add_new_sign, add_r_o, add_exception1, add_exception2, add_exception3, 
        add_exception_o, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [7:0] add_final_exponent;
  input [24:0] add_final_sum;
  output [31:0] add_r_o;
  input clk, reset, new_sign, add_new_sign, add_exception1, add_exception2,
         add_exception3, s;
  output new_sign2, add_exception_o, s2;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N69, N70, N71, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   [31:0] add_r;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[21] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n94), .Q(new_sign2)
         );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n94), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n94), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n93), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n92), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n91), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n90), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n90), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n90), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n90), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n90), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n89), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n89), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n89), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n6), .CLK(clk), .RSTB(n89), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n12), .CLK(clk), .RSTB(n89), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n18), .CLK(clk), .RSTB(n89), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n24), .CLK(clk), .RSTB(n88), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n52), .CLK(clk), .RSTB(n88), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n58), .CLK(clk), .RSTB(n88), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n64), .CLK(clk), .RSTB(n88), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n88), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n88), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n87), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n87), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n87), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n87), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n10), .CLK(clk), .RSTB(n87), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n16), .CLK(clk), .RSTB(n86), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n22), .CLK(clk), .RSTB(n86), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n50), .CLK(clk), .RSTB(n86), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n56), .CLK(clk), .RSTB(n86), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n62), .CLK(clk), .RSTB(n86), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n86), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n86), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n85), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n85), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n85), 
        .Q(new_exponent2[0]) );
  DFFARX1 \add_r_o_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[31]) );
  DFFARX1 \add_r_o_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[30]) );
  DFFARX1 \add_r_o_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[29]) );
  DFFARX1 \add_r_o_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[28]) );
  DFFARX1 \add_r_o_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[27]) );
  DFFARX1 \add_r_o_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[26]) );
  DFFARX1 \add_r_o_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[25]) );
  DFFARX1 \add_r_o_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[24]) );
  DFFARX1 \add_r_o_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n85), .Q(
        add_r_o[23]) );
  DFFARX1 \add_r_o_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[22]) );
  DFFARX1 \add_r_o_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[21]) );
  DFFARX1 \add_r_o_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[20]) );
  DFFARX1 \add_r_o_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[19]) );
  DFFARX1 \add_r_o_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[18]) );
  DFFARX1 \add_r_o_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[17]) );
  DFFARX1 \add_r_o_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[16]) );
  DFFARX1 \add_r_o_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[15]) );
  DFFARX1 \add_r_o_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[14]) );
  DFFARX1 \add_r_o_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[13]) );
  DFFARX1 \add_r_o_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[12]) );
  DFFARX1 \add_r_o_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n84), .Q(
        add_r_o[11]) );
  DFFARX1 \add_r_o_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[10]) );
  DFFARX1 \add_r_o_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[9]) );
  DFFARX1 \add_r_o_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[8]) );
  DFFARX1 \add_r_o_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[7]) );
  DFFARX1 \add_r_o_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[6]) );
  DFFARX1 \add_r_o_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[5]) );
  DFFARX1 \add_r_o_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[4]) );
  DFFARX1 \add_r_o_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[3]) );
  DFFARX1 \add_r_o_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[2]) );
  DFFARX1 \add_r_o_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[1]) );
  DFFARX1 \add_r_o_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n83), .Q(
        add_r_o[0]) );
  DFFARX1 add_exception_o_reg ( .D(n97), .CLK(clk), .RSTB(n83), .Q(
        add_exception_o) );
  AO222X1 U51 ( .IN1(N26), .IN2(n78), .IN3(N77), .IN4(n73), .IN5(
        product_shift[9]), .IN6(n69), .Q(product2[9]) );
  AO222X1 U52 ( .IN1(N25), .IN2(n78), .IN3(N76), .IN4(n73), .IN5(
        product_shift[8]), .IN6(n72), .Q(product2[8]) );
  AO222X1 U53 ( .IN1(N24), .IN2(n78), .IN3(N75), .IN4(n73), .IN5(
        product_shift[7]), .IN6(n72), .Q(product2[7]) );
  AO222X1 U54 ( .IN1(N23), .IN2(n78), .IN3(N74), .IN4(n73), .IN5(
        product_shift[6]), .IN6(n72), .Q(product2[6]) );
  AO222X1 U55 ( .IN1(N22), .IN2(n78), .IN3(N73), .IN4(n73), .IN5(
        product_shift[5]), .IN6(n72), .Q(product2[5]) );
  AO222X1 U56 ( .IN1(N67), .IN2(n78), .IN3(N118), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n72), .Q(product2[50]) );
  AO222X1 U57 ( .IN1(N21), .IN2(n78), .IN3(N72), .IN4(n73), .IN5(
        product_shift[4]), .IN6(n72), .Q(product2[4]) );
  AO222X1 U58 ( .IN1(N66), .IN2(n78), .IN3(N117), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n72), .Q(product2[49]) );
  AO222X1 U59 ( .IN1(N65), .IN2(n78), .IN3(N116), .IN4(n73), .IN5(
        product_shift[48]), .IN6(n72), .Q(product2[48]) );
  AO222X1 U60 ( .IN1(N64), .IN2(n78), .IN3(N115), .IN4(n73), .IN5(
        product_shift[47]), .IN6(n72), .Q(product2[47]) );
  AO222X1 U61 ( .IN1(N63), .IN2(n78), .IN3(N114), .IN4(n73), .IN5(
        product_shift[46]), .IN6(n72), .Q(product2[46]) );
  AO222X1 U62 ( .IN1(N62), .IN2(n78), .IN3(N113), .IN4(n73), .IN5(
        product_shift[45]), .IN6(n72), .Q(product2[45]) );
  AO222X1 U63 ( .IN1(N61), .IN2(n79), .IN3(N112), .IN4(n74), .IN5(
        product_shift[44]), .IN6(n71), .Q(product2[44]) );
  AO222X1 U64 ( .IN1(N60), .IN2(n79), .IN3(N111), .IN4(n74), .IN5(
        product_shift[43]), .IN6(n71), .Q(product2[43]) );
  AO222X1 U65 ( .IN1(N59), .IN2(n79), .IN3(N110), .IN4(n74), .IN5(
        product_shift[42]), .IN6(n71), .Q(product2[42]) );
  AO222X1 U66 ( .IN1(N58), .IN2(n79), .IN3(N109), .IN4(n74), .IN5(
        product_shift[41]), .IN6(n71), .Q(product2[41]) );
  AO222X1 U67 ( .IN1(N57), .IN2(n79), .IN3(N108), .IN4(n74), .IN5(
        product_shift[40]), .IN6(n71), .Q(product2[40]) );
  AO222X1 U68 ( .IN1(N20), .IN2(n79), .IN3(N71), .IN4(n74), .IN5(
        product_shift[3]), .IN6(n71), .Q(product2[3]) );
  AO222X1 U69 ( .IN1(N56), .IN2(n79), .IN3(N107), .IN4(n74), .IN5(
        product_shift[39]), .IN6(n71), .Q(product2[39]) );
  AO222X1 U70 ( .IN1(N55), .IN2(n79), .IN3(N106), .IN4(n74), .IN5(
        product_shift[38]), .IN6(n71), .Q(product2[38]) );
  AO222X1 U71 ( .IN1(N54), .IN2(n79), .IN3(N105), .IN4(n74), .IN5(
        product_shift[37]), .IN6(n71), .Q(product2[37]) );
  AO222X1 U72 ( .IN1(N53), .IN2(n79), .IN3(N104), .IN4(n74), .IN5(
        product_shift[36]), .IN6(n71), .Q(product2[36]) );
  AO222X1 U73 ( .IN1(N52), .IN2(n79), .IN3(N103), .IN4(n74), .IN5(
        product_shift[35]), .IN6(n71), .Q(product2[35]) );
  AO222X1 U74 ( .IN1(N51), .IN2(n79), .IN3(N102), .IN4(n74), .IN5(
        product_shift[34]), .IN6(n71), .Q(product2[34]) );
  AO222X1 U75 ( .IN1(N50), .IN2(n80), .IN3(N101), .IN4(n75), .IN5(n8), .IN6(
        n71), .Q(product2[33]) );
  AO222X1 U76 ( .IN1(N49), .IN2(n80), .IN3(N100), .IN4(n75), .IN5(n14), .IN6(
        n70), .Q(product2[32]) );
  AO222X1 U77 ( .IN1(N48), .IN2(n80), .IN3(N99), .IN4(n75), .IN5(n20), .IN6(
        n70), .Q(product2[31]) );
  AO222X1 U78 ( .IN1(N47), .IN2(n80), .IN3(N98), .IN4(n75), .IN5(n26), .IN6(
        n70), .Q(product2[30]) );
  AO222X1 U79 ( .IN1(N19), .IN2(n80), .IN3(N70), .IN4(n75), .IN5(
        product_shift[2]), .IN6(n70), .Q(product2[2]) );
  AO222X1 U80 ( .IN1(N46), .IN2(n80), .IN3(N97), .IN4(n75), .IN5(n54), .IN6(
        n70), .Q(product2[29]) );
  AO222X1 U81 ( .IN1(N45), .IN2(n80), .IN3(N96), .IN4(n75), .IN5(n60), .IN6(
        n70), .Q(product2[28]) );
  AO222X1 U82 ( .IN1(N44), .IN2(n80), .IN3(N95), .IN4(n75), .IN5(n66), .IN6(
        n70), .Q(product2[27]) );
  AO222X1 U83 ( .IN1(N43), .IN2(n80), .IN3(N94), .IN4(n75), .IN5(n68), .IN6(
        n70), .Q(product2[26]) );
  AO222X1 U84 ( .IN1(N42), .IN2(n80), .IN3(N93), .IN4(n75), .IN5(
        product_shift[25]), .IN6(n70), .Q(product2[25]) );
  AO222X1 U85 ( .IN1(N41), .IN2(n80), .IN3(N92), .IN4(n75), .IN5(
        product_shift[24]), .IN6(n70), .Q(product2[24]) );
  AO222X1 U86 ( .IN1(N40), .IN2(n80), .IN3(N91), .IN4(n75), .IN5(
        product_shift[23]), .IN6(n70), .Q(product2[23]) );
  AO222X1 U87 ( .IN1(N39), .IN2(n81), .IN3(N90), .IN4(n76), .IN5(
        product_shift[22]), .IN6(n70), .Q(product2[22]) );
  AO222X1 U89 ( .IN1(N37), .IN2(n81), .IN3(N88), .IN4(n76), .IN5(
        product_shift[20]), .IN6(n69), .Q(product2[20]) );
  AO222X1 U90 ( .IN1(N18), .IN2(n81), .IN3(N69), .IN4(n76), .IN5(n69), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U91 ( .IN1(N36), .IN2(n81), .IN3(N87), .IN4(n76), .IN5(
        product_shift[19]), .IN6(n69), .Q(product2[19]) );
  AO222X1 U92 ( .IN1(N35), .IN2(n81), .IN3(N86), .IN4(n76), .IN5(
        product_shift[18]), .IN6(n69), .Q(product2[18]) );
  AO222X1 U93 ( .IN1(N34), .IN2(n81), .IN3(N85), .IN4(n76), .IN5(
        product_shift[17]), .IN6(n69), .Q(product2[17]) );
  AO222X1 U94 ( .IN1(N33), .IN2(n81), .IN3(N84), .IN4(n76), .IN5(
        product_shift[16]), .IN6(n69), .Q(product2[16]) );
  AO222X1 U95 ( .IN1(N32), .IN2(n81), .IN3(N83), .IN4(n76), .IN5(
        product_shift[15]), .IN6(n69), .Q(product2[15]) );
  AO222X1 U96 ( .IN1(N31), .IN2(n81), .IN3(N82), .IN4(n76), .IN5(
        product_shift[14]), .IN6(n69), .Q(product2[14]) );
  AO222X1 U97 ( .IN1(N30), .IN2(n81), .IN3(N81), .IN4(n76), .IN5(
        product_shift[13]), .IN6(n69), .Q(product2[13]) );
  AO222X1 U98 ( .IN1(N29), .IN2(n81), .IN3(N80), .IN4(n76), .IN5(
        product_shift[12]), .IN6(n69), .Q(product2[12]) );
  AO222X1 U99 ( .IN1(N28), .IN2(n82), .IN3(N79), .IN4(n77), .IN5(
        product_shift[11]), .IN6(n69), .Q(product2[11]) );
  AO222X1 U100 ( .IN1(N27), .IN2(n82), .IN3(N78), .IN4(n77), .IN5(
        product_shift[10]), .IN6(n70), .Q(product2[10]) );
  XNOR2X1 U102 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n29) );
  AND2X1 U103 ( .IN1(product_shift[1]), .IN2(n95), .Q(n28) );
  AND2X1 U104 ( .IN1(n30), .IN2(add_final_sum[6]), .Q(add_r[6]) );
  AND2X1 U105 ( .IN1(n30), .IN2(add_final_sum[5]), .Q(add_r[5]) );
  AND2X1 U106 ( .IN1(n30), .IN2(add_final_sum[4]), .Q(add_r[4]) );
  AND2X1 U107 ( .IN1(add_new_sign), .IN2(n30), .Q(add_r[31]) );
  AND2X1 U108 ( .IN1(n30), .IN2(add_final_sum[21]), .Q(add_r[21]) );
  AND2X1 U109 ( .IN1(n30), .IN2(add_final_sum[20]), .Q(add_r[20]) );
  AND2X1 U110 ( .IN1(n30), .IN2(add_final_sum[1]), .Q(add_r[1]) );
  AND2X1 U111 ( .IN1(n30), .IN2(add_final_sum[16]), .Q(add_r[16]) );
  AND2X1 U112 ( .IN1(n30), .IN2(add_final_sum[15]), .Q(add_r[15]) );
  AND2X1 U113 ( .IN1(n30), .IN2(add_final_sum[14]), .Q(add_r[14]) );
  AND2X1 U114 ( .IN1(n30), .IN2(add_final_sum[13]), .Q(add_r[13]) );
  AND2X1 U115 ( .IN1(n30), .IN2(add_final_sum[12]), .Q(add_r[12]) );
  AND2X1 U116 ( .IN1(n30), .IN2(add_final_sum[11]), .Q(add_r[11]) );
  OR4X1 U117 ( .IN1(n97), .IN2(n34), .IN3(add_final_sum[24]), .IN4(
        add_final_sum[23]), .Q(n32) );
  OA221X1 U118 ( .IN1(n35), .IN2(n36), .IN3(n37), .IN4(n38), .IN5(n39), .Q(n33) );
  NOR3X0 U119 ( .IN1(add_exception1), .IN2(add_exception3), .IN3(
        add_exception2), .QN(n39) );
  NAND4X0 U120 ( .IN1(add_final_exponent[7]), .IN2(add_final_exponent[6]), 
        .IN3(add_final_exponent[5]), .IN4(add_final_exponent[4]), .QN(n38) );
  NAND4X0 U121 ( .IN1(add_final_exponent[3]), .IN2(add_final_exponent[2]), 
        .IN3(add_final_exponent[1]), .IN4(add_final_exponent[0]), .QN(n37) );
  NAND4X0 U122 ( .IN1(n34), .IN2(n116), .IN3(n115), .IN4(n114), .QN(n36) );
  NAND4X0 U123 ( .IN1(n40), .IN2(n41), .IN3(n42), .IN4(n43), .QN(n34) );
  NOR4X0 U124 ( .IN1(n44), .IN2(add_final_sum[4]), .IN3(add_final_sum[6]), 
        .IN4(add_final_sum[5]), .QN(n43) );
  NAND3X0 U125 ( .IN1(n104), .IN2(n103), .IN3(n105), .QN(n44) );
  NOR4X0 U126 ( .IN1(n45), .IN2(add_final_sum[1]), .IN3(add_final_sum[21]), 
        .IN4(add_final_sum[20]), .QN(n42) );
  NAND3X0 U127 ( .IN1(n107), .IN2(n106), .IN3(n98), .QN(n45) );
  NOR4X0 U128 ( .IN1(n46), .IN2(add_final_sum[14]), .IN3(add_final_sum[16]), 
        .IN4(add_final_sum[15]), .QN(n41) );
  NAND3X0 U129 ( .IN1(n100), .IN2(n99), .IN3(n101), .QN(n46) );
  NOR4X0 U130 ( .IN1(n47), .IN2(add_final_sum[11]), .IN3(add_final_sum[13]), 
        .IN4(add_final_sum[12]), .QN(n40) );
  NAND4X0 U131 ( .IN1(n113), .IN2(n112), .IN3(n48), .IN4(n111), .QN(n35) );
  booth5_DW01_add_0 add_91 ( .A({product_shift[49], product_shift[49:34], n8, 
        n14, n20, n26, n54, n60, n66, n68, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n10, n16, n22, n50, n56, n62, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N118, N117, 
        N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, 
        N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, 
        N91, N90, SYNOPSYS_UNCONNECTED__0, N88, N87, N86, N85, N84, N83, N82, 
        N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth5_DW01_add_1 add_84 ( .A({product_shift[49], product_shift[49:34], n8, 
        n14, n20, n26, n54, n60, n66, n68, product_shift[25:0]}), .B({
        combined_b[24:8], n6, n12, n18, n24, n52, n58, n64, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, SYNOPSYS_UNCONNECTED__2, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U7 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U8 ( .INP(n5), .ZN(n6) );
  INVX0 U9 ( .INP(product_shift[33]), .ZN(n7) );
  INVX0 U10 ( .INP(n7), .ZN(n8) );
  INVX0 U11 ( .INP(combined_negative_b[6]), .ZN(n9) );
  INVX0 U12 ( .INP(n9), .ZN(n10) );
  INVX0 U13 ( .INP(combined_b[6]), .ZN(n11) );
  INVX0 U14 ( .INP(n11), .ZN(n12) );
  INVX0 U15 ( .INP(product_shift[32]), .ZN(n13) );
  INVX0 U16 ( .INP(n13), .ZN(n14) );
  INVX0 U17 ( .INP(combined_negative_b[5]), .ZN(n15) );
  INVX0 U18 ( .INP(n15), .ZN(n16) );
  INVX0 U19 ( .INP(combined_b[5]), .ZN(n17) );
  INVX0 U20 ( .INP(n17), .ZN(n18) );
  INVX0 U21 ( .INP(product_shift[31]), .ZN(n19) );
  INVX0 U22 ( .INP(n19), .ZN(n20) );
  INVX0 U23 ( .INP(combined_negative_b[4]), .ZN(n21) );
  INVX0 U24 ( .INP(n21), .ZN(n22) );
  INVX0 U25 ( .INP(combined_b[4]), .ZN(n23) );
  INVX0 U26 ( .INP(n23), .ZN(n24) );
  INVX0 U27 ( .INP(product_shift[30]), .ZN(n25) );
  INVX0 U28 ( .INP(n25), .ZN(n26) );
  INVX0 U29 ( .INP(combined_negative_b[3]), .ZN(n49) );
  INVX0 U30 ( .INP(n49), .ZN(n50) );
  INVX0 U31 ( .INP(combined_b[3]), .ZN(n51) );
  INVX0 U32 ( .INP(n51), .ZN(n52) );
  INVX0 U33 ( .INP(product_shift[29]), .ZN(n53) );
  INVX0 U34 ( .INP(n53), .ZN(n54) );
  INVX0 U35 ( .INP(combined_negative_b[2]), .ZN(n55) );
  INVX0 U36 ( .INP(n55), .ZN(n56) );
  INVX0 U37 ( .INP(combined_b[2]), .ZN(n57) );
  INVX0 U38 ( .INP(n57), .ZN(n58) );
  INVX0 U39 ( .INP(product_shift[28]), .ZN(n59) );
  INVX0 U40 ( .INP(n59), .ZN(n60) );
  INVX0 U41 ( .INP(combined_negative_b[1]), .ZN(n61) );
  INVX0 U42 ( .INP(n61), .ZN(n62) );
  INVX0 U43 ( .INP(combined_b[1]), .ZN(n63) );
  INVX0 U44 ( .INP(n63), .ZN(n64) );
  INVX0 U45 ( .INP(n30), .ZN(n96) );
  NAND2X1 U46 ( .IN1(n32), .IN2(n33), .QN(n31) );
  NAND2X1 U47 ( .IN1(n32), .IN2(n31), .QN(n30) );
  NBUFFX2 U48 ( .INP(n27), .Z(n80) );
  NBUFFX2 U49 ( .INP(n27), .Z(n79) );
  NBUFFX2 U50 ( .INP(n27), .Z(n78) );
  NBUFFX2 U88 ( .INP(n27), .Z(n81) );
  NOR2X0 U101 ( .IN1(n96), .IN2(n108), .QN(add_r[0]) );
  NOR2X0 U132 ( .IN1(n96), .IN2(n107), .QN(add_r[2]) );
  NOR2X0 U133 ( .IN1(n96), .IN2(n106), .QN(add_r[3]) );
  NOR2X0 U134 ( .IN1(n96), .IN2(n105), .QN(add_r[7]) );
  NOR2X0 U135 ( .IN1(n96), .IN2(n104), .QN(add_r[8]) );
  NOR2X0 U136 ( .IN1(n96), .IN2(n103), .QN(add_r[9]) );
  NOR2X0 U137 ( .IN1(n96), .IN2(n102), .QN(add_r[10]) );
  NOR2X0 U138 ( .IN1(n96), .IN2(n101), .QN(add_r[17]) );
  NOR2X0 U139 ( .IN1(n96), .IN2(n100), .QN(add_r[18]) );
  NOR2X0 U140 ( .IN1(n96), .IN2(n99), .QN(add_r[19]) );
  NOR2X0 U141 ( .IN1(n96), .IN2(n98), .QN(add_r[22]) );
  NOR2X0 U142 ( .IN1(n116), .IN2(n31), .QN(add_r[23]) );
  NOR2X0 U143 ( .IN1(n115), .IN2(n31), .QN(add_r[24]) );
  NOR2X0 U144 ( .IN1(n114), .IN2(n31), .QN(add_r[25]) );
  NOR2X0 U145 ( .IN1(n113), .IN2(n31), .QN(add_r[26]) );
  NOR2X0 U146 ( .IN1(n112), .IN2(n31), .QN(add_r[27]) );
  NOR2X0 U147 ( .IN1(n111), .IN2(n31), .QN(add_r[28]) );
  NBUFFX2 U148 ( .INP(n27), .Z(n82) );
  INVX0 U149 ( .INP(n33), .ZN(n97) );
  NBUFFX2 U150 ( .INP(n29), .Z(n70) );
  NBUFFX2 U151 ( .INP(n29), .Z(n71) );
  NBUFFX2 U152 ( .INP(n29), .Z(n69) );
  NBUFFX2 U153 ( .INP(n29), .Z(n72) );
  NBUFFX2 U154 ( .INP(n28), .Z(n75) );
  NBUFFX2 U155 ( .INP(n28), .Z(n74) );
  NBUFFX2 U156 ( .INP(n28), .Z(n73) );
  NBUFFX2 U157 ( .INP(n28), .Z(n76) );
  NBUFFX2 U158 ( .INP(n28), .Z(n77) );
  NBUFFX2 U159 ( .INP(reset), .Z(n83) );
  NBUFFX2 U160 ( .INP(reset), .Z(n84) );
  NBUFFX2 U161 ( .INP(reset), .Z(n85) );
  NBUFFX2 U162 ( .INP(reset), .Z(n86) );
  NBUFFX2 U163 ( .INP(reset), .Z(n87) );
  NBUFFX2 U164 ( .INP(reset), .Z(n88) );
  NBUFFX2 U165 ( .INP(reset), .Z(n89) );
  NBUFFX2 U166 ( .INP(reset), .Z(n90) );
  NBUFFX2 U167 ( .INP(reset), .Z(n91) );
  NBUFFX2 U168 ( .INP(reset), .Z(n93) );
  NBUFFX2 U169 ( .INP(reset), .Z(n94) );
  NBUFFX2 U170 ( .INP(reset), .Z(n92) );
  NOR2X0 U171 ( .IN1(n95), .IN2(product_shift[1]), .QN(n27) );
  NOR2X0 U172 ( .IN1(n110), .IN2(n31), .QN(add_r[29]) );
  INVX0 U173 ( .INP(add_final_exponent[6]), .ZN(n110) );
  NOR2X0 U174 ( .IN1(n109), .IN2(n31), .QN(add_r[30]) );
  INVX0 U175 ( .INP(add_final_exponent[7]), .ZN(n109) );
  INVX0 U176 ( .INP(add_final_sum[10]), .ZN(n102) );
  INVX0 U177 ( .INP(add_final_sum[0]), .ZN(n108) );
  NOR2X0 U178 ( .IN1(add_final_exponent[7]), .IN2(add_final_exponent[6]), .QN(
        n48) );
  NAND2X1 U179 ( .IN1(n108), .IN2(n102), .QN(n47) );
  INVX0 U180 ( .INP(add_final_exponent[2]), .ZN(n114) );
  INVX0 U181 ( .INP(add_final_exponent[5]), .ZN(n111) );
  INVX0 U182 ( .INP(add_final_exponent[1]), .ZN(n115) );
  INVX0 U183 ( .INP(add_final_exponent[4]), .ZN(n112) );
  INVX0 U184 ( .INP(add_final_exponent[0]), .ZN(n116) );
  INVX0 U185 ( .INP(add_final_exponent[3]), .ZN(n113) );
  INVX0 U186 ( .INP(add_final_sum[7]), .ZN(n105) );
  INVX0 U187 ( .INP(add_final_sum[22]), .ZN(n98) );
  INVX0 U188 ( .INP(add_final_sum[17]), .ZN(n101) );
  INVX0 U189 ( .INP(add_final_sum[9]), .ZN(n103) );
  INVX0 U190 ( .INP(add_final_sum[3]), .ZN(n106) );
  INVX0 U191 ( .INP(add_final_sum[19]), .ZN(n99) );
  INVX0 U192 ( .INP(add_final_sum[8]), .ZN(n104) );
  INVX0 U193 ( .INP(add_final_sum[2]), .ZN(n107) );
  INVX0 U194 ( .INP(add_final_sum[18]), .ZN(n100) );
  INVX0 U195 ( .INP(product_shift[0]), .ZN(n95) );
  INVX0 U197 ( .INP(product_shift[27]), .ZN(n65) );
  INVX0 U198 ( .INP(n65), .ZN(n66) );
  INVX0 U199 ( .INP(product_shift[26]), .ZN(n67) );
  INVX0 U200 ( .INP(n67), .ZN(n68) );
endmodule


module booth6_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X1 U2 ( .IN1(A[46]), .IN2(carry[46]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[46]), .IN2(carry[46]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[46]), .IN2(A[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[47]) );
  XOR3X1 U6 ( .IN1(carry[47]), .IN2(B[47]), .IN3(A[47]), .Q(SUM[47]) );
  NAND2X0 U7 ( .IN1(A[47]), .IN2(carry[47]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[47]), .IN2(carry[47]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[47]), .IN2(A[47]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[48]) );
  XOR3X2 U11 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U12 ( .IN1(A[48]), .IN2(B[48]), .QN(n7) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(carry[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(B[48]), .IN2(carry[48]), .QN(n9) );
  NAND3X0 U15 ( .IN1(n7), .IN2(n8), .IN3(n9), .QN(carry[49]) );
  XOR2X1 U16 ( .IN1(A[49]), .IN2(B[49]), .Q(n10) );
  XOR2X1 U17 ( .IN1(n10), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U18 ( .IN1(A[49]), .IN2(B[49]), .QN(n11) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(carry[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(B[49]), .IN2(carry[49]), .QN(n13) );
  NAND3X0 U21 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[50]) );
  DELLN2X2 U22 ( .INP(carry[45]), .Z(n14) );
  NAND2X0 U23 ( .IN1(n25), .IN2(B[27]), .QN(n23) );
  XOR3X2 U24 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U25 ( .IN1(A[44]), .IN2(B[44]), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[44]), .IN2(carry[44]), .QN(n16) );
  NAND2X0 U27 ( .IN1(B[44]), .IN2(carry[44]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n16), .IN2(n17), .IN3(n15), .QN(carry[45]) );
  XOR2X1 U29 ( .IN1(A[45]), .IN2(B[45]), .Q(n18) );
  XOR2X1 U30 ( .IN1(n18), .IN2(n14), .Q(SUM[45]) );
  NAND2X0 U31 ( .IN1(A[45]), .IN2(B[45]), .QN(n19) );
  NAND2X0 U32 ( .IN1(A[45]), .IN2(carry[45]), .QN(n20) );
  NAND2X0 U33 ( .IN1(B[45]), .IN2(carry[45]), .QN(n21) );
  NAND3X0 U34 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[46]) );
  XOR3X1 U35 ( .IN1(B[27]), .IN2(n25), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U36 ( .IN1(A[27]), .IN2(B[27]), .QN(n22) );
  NAND2X0 U37 ( .IN1(n25), .IN2(A[27]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n24), .IN3(n23), .QN(carry[28]) );
  AND2X4 U39 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  XOR2X1 U40 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_35 ( .A(n12), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  XOR3X1 U1 ( .IN1(carry[43]), .IN2(B[43]), .IN3(A[43]), .Q(SUM[43]) );
  NAND2X1 U2 ( .IN1(A[43]), .IN2(carry[43]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[43]), .IN2(carry[43]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[43]), .IN2(A[43]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[44]) );
  XOR3X2 U6 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U7 ( .IN1(A[38]), .IN2(B[38]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[38]), .IN2(carry[38]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[38]), .IN2(carry[38]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[39]) );
  XOR2X1 U11 ( .IN1(A[39]), .IN2(B[39]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U13 ( .IN1(A[39]), .IN2(B[39]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[39]), .IN2(carry[39]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[39]), .IN2(carry[39]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[40]) );
  INVX0 U17 ( .INP(A[35]), .ZN(n11) );
  INVX0 U18 ( .INP(n11), .ZN(n12) );
  NAND2X0 U19 ( .IN1(n24), .IN2(B[27]), .QN(n22) );
  DELLN2X2 U20 ( .INP(carry[41]), .Z(n13) );
  XOR3X2 U21 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  NAND2X0 U22 ( .IN1(A[40]), .IN2(B[40]), .QN(n14) );
  NAND2X0 U23 ( .IN1(A[40]), .IN2(carry[40]), .QN(n15) );
  NAND2X0 U24 ( .IN1(B[40]), .IN2(carry[40]), .QN(n16) );
  NAND3X0 U25 ( .IN1(n16), .IN2(n15), .IN3(n14), .QN(carry[41]) );
  XOR2X1 U26 ( .IN1(A[41]), .IN2(B[41]), .Q(n17) );
  XOR2X1 U27 ( .IN1(n17), .IN2(n13), .Q(SUM[41]) );
  NAND2X0 U28 ( .IN1(A[41]), .IN2(B[41]), .QN(n18) );
  NAND2X0 U29 ( .IN1(A[41]), .IN2(carry[41]), .QN(n19) );
  NAND2X0 U30 ( .IN1(B[41]), .IN2(carry[41]), .QN(n20) );
  NAND3X0 U31 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[42]) );
  XOR3X1 U32 ( .IN1(B[27]), .IN2(n24), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U33 ( .IN1(A[27]), .IN2(B[27]), .QN(n21) );
  NAND2X0 U34 ( .IN1(n24), .IN2(A[27]), .QN(n23) );
  NAND3X0 U35 ( .IN1(n21), .IN2(n23), .IN3(n22), .QN(carry[28]) );
  AND2X4 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(n24) );
  XOR2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_0 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n6, n7, n8, n3, n4, n5, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[20] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n71), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n71), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(n4), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(n9), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n15), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n21), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n27), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n33), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n39), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n45), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n64), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n11), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n17), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n23), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n29), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n35), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n41), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n47), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n62), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n60), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n60), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n60), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n60), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n60), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n60), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n60), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n60), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n60), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n60), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n56), .IN3(N75), .IN4(n7), .IN5(
        product_shift[9]), .IN6(n8), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n56), .IN3(N74), .IN4(n7), .IN5(
        product_shift[8]), .IN6(n8), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n56), .IN3(N73), .IN4(n7), .IN5(
        product_shift[7]), .IN6(n8), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n56), .IN3(N72), .IN4(n7), .IN5(
        product_shift[6]), .IN6(n8), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n56), .IN3(N71), .IN4(n7), .IN5(
        product_shift[5]), .IN6(n8), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(n56), .IN2(N65), .IN3(N116), .IN4(n7), .IN5(
        product_shift[49]), .IN6(n8), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n56), .IN3(N70), .IN4(n7), .IN5(
        product_shift[4]), .IN6(n8), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n56), .IN3(N115), .IN4(n7), .IN5(
        product_shift[49]), .IN6(n8), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n56), .IN3(N114), .IN4(n7), .IN5(
        product_shift[48]), .IN6(n8), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n56), .IN3(N113), .IN4(n7), .IN5(
        product_shift[47]), .IN6(n53), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n56), .IN3(N112), .IN4(n7), .IN5(
        product_shift[46]), .IN6(n53), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n56), .IN3(N111), .IN4(n55), .IN5(
        product_shift[45]), .IN6(n52), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n57), .IN3(N110), .IN4(n54), .IN5(
        product_shift[44]), .IN6(n53), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n57), .IN3(N109), .IN4(n54), .IN5(
        product_shift[43]), .IN6(n53), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n57), .IN3(N108), .IN4(n54), .IN5(
        product_shift[42]), .IN6(n53), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n57), .IN3(N107), .IN4(n54), .IN5(
        product_shift[41]), .IN6(n53), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n57), .IN3(N106), .IN4(n54), .IN5(
        product_shift[40]), .IN6(n53), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n57), .IN3(N69), .IN4(n54), .IN5(
        product_shift[3]), .IN6(n53), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n57), .IN3(N105), .IN4(n54), .IN5(
        product_shift[39]), .IN6(n53), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n57), .IN3(N104), .IN4(n54), .IN5(
        product_shift[38]), .IN6(n53), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n57), .IN3(N103), .IN4(n54), .IN5(
        product_shift[37]), .IN6(n53), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n57), .IN3(N102), .IN4(n54), .IN5(
        product_shift[36]), .IN6(n53), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n57), .IN3(N101), .IN4(n54), .IN5(
        product_shift[35]), .IN6(n53), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n57), .IN3(N100), .IN4(n54), .IN5(n13), .IN6(
        n53), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n58), .IN3(N99), .IN4(n55), .IN5(n19), .IN6(
        n53), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n58), .IN3(N98), .IN4(n55), .IN5(n25), .IN6(
        n52), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n58), .IN3(N97), .IN4(n55), .IN5(n31), .IN6(
        n52), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n58), .IN3(N96), .IN4(n55), .IN5(n37), .IN6(
        n52), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n58), .IN3(N68), .IN4(n55), .IN5(
        product_shift[2]), .IN6(n52), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n58), .IN3(N95), .IN4(n55), .IN5(n43), .IN6(
        n52), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n58), .IN3(N94), .IN4(n55), .IN5(n49), .IN6(
        n52), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n58), .IN3(N93), .IN4(n55), .IN5(n51), .IN6(
        n52), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n58), .IN3(N92), .IN4(n55), .IN5(
        product_shift[26]), .IN6(n52), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n58), .IN3(N91), .IN4(n55), .IN5(
        product_shift[25]), .IN6(n52), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n58), .IN3(N90), .IN4(n55), .IN5(
        product_shift[24]), .IN6(n52), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n58), .IN3(N89), .IN4(n55), .IN5(
        product_shift[23]), .IN6(n52), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n59), .IN3(N88), .IN4(n7), .IN5(
        product_shift[22]), .IN6(n52), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n59), .IN3(N87), .IN4(n7), .IN5(
        product_shift[21]), .IN6(n8), .Q(product2[21]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n59), .IN3(N67), .IN4(n55), .IN5(n8), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n59), .IN3(N85), .IN4(n7), .IN5(
        product_shift[19]), .IN6(n8), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n59), .IN3(N84), .IN4(n7), .IN5(
        product_shift[18]), .IN6(n8), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n59), .IN3(N83), .IN4(n7), .IN5(
        product_shift[17]), .IN6(n8), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n59), .IN3(N82), .IN4(n7), .IN5(
        product_shift[16]), .IN6(n8), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n59), .IN3(N81), .IN4(n7), .IN5(
        product_shift[15]), .IN6(n8), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n59), .IN3(N80), .IN4(n7), .IN5(
        product_shift[14]), .IN6(n8), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n59), .IN3(N79), .IN4(n7), .IN5(
        product_shift[13]), .IN6(n8), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n59), .IN3(N78), .IN4(n7), .IN5(
        product_shift[12]), .IN6(n8), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n59), .IN3(N77), .IN4(n54), .IN5(
        product_shift[11]), .IN6(n52), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n59), .IN3(N76), .IN4(n54), .IN5(
        product_shift[10]), .IN6(n52), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n8) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n72), .Q(n7) );
  booth6_0_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:35], 
        n13, n19, n25, n31, n37, n43, n49, n51, product_shift[26:0]}), .B({
        combined_negative_b[24:9], n11, n17, n23, n29, n35, n41, n47, 
        combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, SYNOPSYS_UNCONNECTED__0, N85, N84, N83, N82, N81, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_0_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:35], 
        n13, n19, n25, n31, n37, n43, n49, n51, product_shift[26:0]}), .B({
        combined_b[24:10], n4, n9, n15, n21, n27, n33, n39, n45, 
        combined_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        SYNOPSYS_UNCONNECTED__2, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, 
        SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_b[9]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  NBUFFX2 U45 ( .INP(reset), .Z(n60) );
  NBUFFX2 U57 ( .INP(reset), .Z(n61) );
  NBUFFX2 U60 ( .INP(reset), .Z(n62) );
  NBUFFX2 U61 ( .INP(reset), .Z(n63) );
  NBUFFX2 U62 ( .INP(reset), .Z(n64) );
  NBUFFX2 U63 ( .INP(reset), .Z(n65) );
  NBUFFX2 U64 ( .INP(reset), .Z(n66) );
  NBUFFX2 U65 ( .INP(reset), .Z(n67) );
  NBUFFX2 U66 ( .INP(reset), .Z(n68) );
  INVX0 U67 ( .INP(combined_b[8]), .ZN(n5) );
  INVX0 U68 ( .INP(n5), .ZN(n9) );
  INVX0 U69 ( .INP(combined_negative_b[8]), .ZN(n10) );
  INVX0 U70 ( .INP(n10), .ZN(n11) );
  INVX0 U71 ( .INP(product_shift[34]), .ZN(n12) );
  INVX0 U72 ( .INP(n12), .ZN(n13) );
  INVX0 U73 ( .INP(combined_b[7]), .ZN(n14) );
  INVX0 U74 ( .INP(n14), .ZN(n15) );
  INVX0 U75 ( .INP(combined_negative_b[7]), .ZN(n16) );
  INVX0 U76 ( .INP(n16), .ZN(n17) );
  INVX0 U77 ( .INP(product_shift[33]), .ZN(n18) );
  INVX0 U78 ( .INP(n18), .ZN(n19) );
  INVX0 U79 ( .INP(combined_b[6]), .ZN(n20) );
  INVX0 U80 ( .INP(n20), .ZN(n21) );
  INVX0 U81 ( .INP(combined_negative_b[6]), .ZN(n22) );
  INVX0 U82 ( .INP(n22), .ZN(n23) );
  INVX0 U83 ( .INP(product_shift[32]), .ZN(n24) );
  INVX0 U84 ( .INP(n24), .ZN(n25) );
  INVX0 U85 ( .INP(combined_b[5]), .ZN(n26) );
  INVX0 U86 ( .INP(n26), .ZN(n27) );
  INVX0 U87 ( .INP(combined_negative_b[5]), .ZN(n28) );
  INVX0 U88 ( .INP(n28), .ZN(n29) );
  INVX0 U89 ( .INP(product_shift[31]), .ZN(n30) );
  INVX0 U90 ( .INP(n30), .ZN(n31) );
  INVX0 U91 ( .INP(combined_b[4]), .ZN(n32) );
  INVX0 U92 ( .INP(n32), .ZN(n33) );
  INVX0 U93 ( .INP(combined_negative_b[4]), .ZN(n34) );
  INVX0 U94 ( .INP(n34), .ZN(n35) );
  INVX0 U95 ( .INP(product_shift[30]), .ZN(n36) );
  INVX0 U96 ( .INP(n36), .ZN(n37) );
  INVX0 U97 ( .INP(combined_b[3]), .ZN(n38) );
  INVX0 U98 ( .INP(n38), .ZN(n39) );
  INVX0 U99 ( .INP(combined_negative_b[3]), .ZN(n40) );
  INVX0 U100 ( .INP(n40), .ZN(n41) );
  INVX0 U101 ( .INP(product_shift[29]), .ZN(n42) );
  INVX0 U102 ( .INP(n42), .ZN(n43) );
  INVX0 U103 ( .INP(combined_b[2]), .ZN(n44) );
  INVX0 U104 ( .INP(n44), .ZN(n45) );
  INVX0 U105 ( .INP(combined_negative_b[2]), .ZN(n46) );
  INVX0 U106 ( .INP(n46), .ZN(n47) );
  INVX0 U107 ( .INP(product_shift[28]), .ZN(n48) );
  INVX0 U108 ( .INP(n48), .ZN(n49) );
  NBUFFX2 U109 ( .INP(n6), .Z(n58) );
  NBUFFX2 U110 ( .INP(n6), .Z(n57) );
  NBUFFX2 U111 ( .INP(n6), .Z(n56) );
  NBUFFX2 U112 ( .INP(n6), .Z(n59) );
  NBUFFX2 U113 ( .INP(n8), .Z(n52) );
  NBUFFX2 U114 ( .INP(n8), .Z(n53) );
  NBUFFX2 U115 ( .INP(n7), .Z(n55) );
  NBUFFX2 U116 ( .INP(n7), .Z(n54) );
  NBUFFX2 U117 ( .INP(reset), .Z(n70) );
  NBUFFX2 U118 ( .INP(reset), .Z(n71) );
  NBUFFX2 U119 ( .INP(reset), .Z(n69) );
  NOR2X0 U120 ( .IN1(n72), .IN2(product_shift[1]), .QN(n6) );
  INVX0 U121 ( .INP(product_shift[0]), .ZN(n72) );
  INVX0 U123 ( .INP(product_shift[27]), .ZN(n50) );
  INVX0 U124 ( .INP(n50), .ZN(n51) );
endmodule


module booth6_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  XOR3X1 U1 ( .IN1(carry[47]), .IN2(B[47]), .IN3(A[47]), .Q(SUM[47]) );
  NAND2X0 U2 ( .IN1(A[47]), .IN2(carry[47]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[47]), .IN2(carry[47]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[47]), .IN2(A[47]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[48]) );
  XOR3X2 U6 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  NAND2X0 U7 ( .IN1(A[40]), .IN2(B[40]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[40]), .IN2(carry[40]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[40]), .IN2(carry[40]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[41]) );
  XOR2X1 U11 ( .IN1(A[41]), .IN2(B[41]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[41]), .Q(SUM[41]) );
  NAND2X0 U13 ( .IN1(A[41]), .IN2(B[41]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[41]), .IN2(carry[41]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[41]), .IN2(carry[41]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[42]) );
  XOR3X1 U17 ( .IN1(carry[43]), .IN2(B[43]), .IN3(A[43]), .Q(SUM[43]) );
  NAND2X0 U18 ( .IN1(A[43]), .IN2(carry[43]), .QN(n11) );
  NAND2X0 U19 ( .IN1(B[43]), .IN2(carry[43]), .QN(n12) );
  NAND2X0 U20 ( .IN1(B[43]), .IN2(A[43]), .QN(n13) );
  NAND3X0 U21 ( .IN1(n11), .IN2(n13), .IN3(n12), .QN(carry[44]) );
  NAND2X0 U22 ( .IN1(n25), .IN2(B[27]), .QN(n23) );
  DELLN2X2 U23 ( .INP(carry[45]), .Z(n14) );
  XOR3X2 U24 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U25 ( .IN1(A[44]), .IN2(B[44]), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[44]), .IN2(carry[44]), .QN(n16) );
  NAND2X0 U27 ( .IN1(B[44]), .IN2(carry[44]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[45]) );
  XOR2X1 U29 ( .IN1(A[45]), .IN2(B[45]), .Q(n18) );
  XOR2X1 U30 ( .IN1(n18), .IN2(n14), .Q(SUM[45]) );
  NAND2X0 U31 ( .IN1(A[45]), .IN2(B[45]), .QN(n19) );
  NAND2X0 U32 ( .IN1(A[45]), .IN2(carry[45]), .QN(n20) );
  NAND2X0 U33 ( .IN1(B[45]), .IN2(carry[45]), .QN(n21) );
  NAND3X0 U34 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[46]) );
  XOR3X1 U35 ( .IN1(B[27]), .IN2(n25), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U36 ( .IN1(A[27]), .IN2(B[27]), .QN(n22) );
  NAND2X0 U37 ( .IN1(n25), .IN2(A[27]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n24), .IN3(n23), .QN(carry[28]) );
  AND2X4 U39 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  XOR2X1 U40 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_19_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X1 U1 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U2 ( .IN1(A[46]), .IN2(carry[46]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[46]), .IN2(carry[46]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[46]), .IN2(A[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[47]) );
  XOR3X2 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U7 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U11 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U13 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  XOR3X1 U17 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U18 ( .IN1(A[42]), .IN2(carry[42]), .QN(n11) );
  NAND2X0 U19 ( .IN1(B[42]), .IN2(carry[42]), .QN(n12) );
  NAND2X0 U20 ( .IN1(B[42]), .IN2(A[42]), .QN(n13) );
  NAND3X0 U21 ( .IN1(n11), .IN2(n13), .IN3(n12), .QN(carry[43]) );
  NAND2X0 U22 ( .IN1(n25), .IN2(B[27]), .QN(n23) );
  DELLN2X2 U23 ( .INP(carry[44]), .Z(n14) );
  XOR3X2 U24 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U25 ( .IN1(A[43]), .IN2(B[43]), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[43]), .IN2(carry[43]), .QN(n16) );
  NAND2X0 U27 ( .IN1(B[43]), .IN2(carry[43]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n17), .IN2(n16), .IN3(n15), .QN(carry[44]) );
  XOR2X1 U29 ( .IN1(A[44]), .IN2(B[44]), .Q(n18) );
  XOR2X1 U30 ( .IN1(n18), .IN2(n14), .Q(SUM[44]) );
  NAND2X0 U31 ( .IN1(A[44]), .IN2(B[44]), .QN(n19) );
  NAND2X0 U32 ( .IN1(A[44]), .IN2(carry[44]), .QN(n20) );
  NAND2X0 U33 ( .IN1(B[44]), .IN2(carry[44]), .QN(n21) );
  NAND3X0 U34 ( .IN1(n20), .IN2(n21), .IN3(n19), .QN(carry[45]) );
  XOR3X1 U35 ( .IN1(B[27]), .IN2(n25), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U36 ( .IN1(A[27]), .IN2(B[27]), .QN(n22) );
  NAND2X0 U37 ( .IN1(n25), .IN2(A[27]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n24), .IN3(n23), .QN(carry[28]) );
  AND2X4 U39 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  XOR2X1 U40 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_19 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[19] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n70), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n70), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n67), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(n9), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n15), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n21), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n27), .CLK(clk), .RSTB(n66), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n33), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n39), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n45), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n65), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n64), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n4), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n13), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n19), .CLK(clk), .RSTB(n64), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n25), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n31), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n37), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n43), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n63), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n62), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n60), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n60), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n60), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n60), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n60), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n60), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n60), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n60), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n60), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n60), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n56), .IN3(N75), .IN4(n73), .IN5(
        product_shift[9]), .IN6(n72), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n56), .IN3(N74), .IN4(n73), .IN5(
        product_shift[8]), .IN6(n72), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n56), .IN3(N73), .IN4(n73), .IN5(
        product_shift[7]), .IN6(n72), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n56), .IN3(N72), .IN4(n73), .IN5(
        product_shift[6]), .IN6(n72), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n56), .IN3(N71), .IN4(n73), .IN5(
        product_shift[5]), .IN6(n72), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n56), .IN3(N116), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n72), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n56), .IN3(N70), .IN4(n73), .IN5(
        product_shift[4]), .IN6(n72), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n56), .IN3(N115), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n72), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n56), .IN3(N114), .IN4(n73), .IN5(
        product_shift[48]), .IN6(n72), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n56), .IN3(N113), .IN4(n73), .IN5(
        product_shift[47]), .IN6(n53), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n56), .IN3(N112), .IN4(n73), .IN5(
        product_shift[46]), .IN6(n53), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n56), .IN3(N111), .IN4(n55), .IN5(
        product_shift[45]), .IN6(n52), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n57), .IN3(N110), .IN4(n54), .IN5(
        product_shift[44]), .IN6(n53), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n57), .IN3(N109), .IN4(n54), .IN5(
        product_shift[43]), .IN6(n53), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n57), .IN3(N108), .IN4(n54), .IN5(
        product_shift[42]), .IN6(n53), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n57), .IN3(N107), .IN4(n54), .IN5(
        product_shift[41]), .IN6(n53), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n57), .IN3(N106), .IN4(n54), .IN5(
        product_shift[40]), .IN6(n53), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n57), .IN3(N69), .IN4(n54), .IN5(
        product_shift[3]), .IN6(n53), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n57), .IN3(N105), .IN4(n54), .IN5(
        product_shift[39]), .IN6(n53), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n57), .IN3(N104), .IN4(n54), .IN5(
        product_shift[38]), .IN6(n53), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n57), .IN3(N103), .IN4(n54), .IN5(
        product_shift[37]), .IN6(n53), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n57), .IN3(N102), .IN4(n54), .IN5(
        product_shift[36]), .IN6(n53), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n57), .IN3(N101), .IN4(n54), .IN5(
        product_shift[35]), .IN6(n53), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n57), .IN3(N100), .IN4(n54), .IN5(n11), .IN6(
        n53), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n58), .IN3(N99), .IN4(n55), .IN5(n17), .IN6(
        n53), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n58), .IN3(N98), .IN4(n55), .IN5(n23), .IN6(
        n52), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n58), .IN3(N97), .IN4(n55), .IN5(n29), .IN6(
        n52), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n58), .IN3(N96), .IN4(n55), .IN5(n35), .IN6(
        n52), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n58), .IN3(N68), .IN4(n55), .IN5(
        product_shift[2]), .IN6(n52), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n58), .IN3(N95), .IN4(n55), .IN5(n41), .IN6(
        n52), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n58), .IN3(N94), .IN4(n55), .IN5(n47), .IN6(
        n52), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n58), .IN3(N93), .IN4(n55), .IN5(n49), .IN6(
        n52), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n58), .IN3(N92), .IN4(n55), .IN5(
        product_shift[26]), .IN6(n52), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n58), .IN3(N91), .IN4(n55), .IN5(
        product_shift[25]), .IN6(n52), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n58), .IN3(N90), .IN4(n55), .IN5(
        product_shift[24]), .IN6(n52), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n58), .IN3(N89), .IN4(n55), .IN5(
        product_shift[23]), .IN6(n52), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n59), .IN3(N88), .IN4(n73), .IN5(
        product_shift[22]), .IN6(n52), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n59), .IN3(N87), .IN4(n73), .IN5(
        product_shift[21]), .IN6(n72), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n59), .IN3(N86), .IN4(n73), .IN5(
        product_shift[20]), .IN6(n72), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n59), .IN3(N67), .IN4(n55), .IN5(n72), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n59), .IN3(N84), .IN4(n73), .IN5(
        product_shift[18]), .IN6(n72), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n59), .IN3(N83), .IN4(n73), .IN5(
        product_shift[17]), .IN6(n72), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n59), .IN3(N82), .IN4(n73), .IN5(
        product_shift[16]), .IN6(n72), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n59), .IN3(N81), .IN4(n73), .IN5(
        product_shift[15]), .IN6(n72), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n59), .IN3(N80), .IN4(n73), .IN5(
        product_shift[14]), .IN6(n72), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n59), .IN3(N79), .IN4(n73), .IN5(
        product_shift[13]), .IN6(n72), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n59), .IN3(N78), .IN4(n73), .IN5(
        product_shift[12]), .IN6(n72), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n59), .IN3(N77), .IN4(n54), .IN5(
        product_shift[11]), .IN6(n52), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n59), .IN3(N76), .IN4(n54), .IN5(
        product_shift[10]), .IN6(n52), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n72) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n71), .Q(n73) );
  booth6_19_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:35], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[26:0]}), .B({
        combined_negative_b[24:9], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, SYNOPSYS_UNCONNECTED__0, N84, N83, N82, N81, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_19_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:35], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[26:0]}), .B({
        combined_b[24:9], n9, n15, n21, n27, n33, n39, n45, combined_b[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, SYNOPSYS_UNCONNECTED__2, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[48]) );
  INVX0 U3 ( .INP(combined_negative_b[8]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U47 ( .INP(combined_b[8]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[34]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[7]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[7]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[33]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[6]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[6]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[32]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[5]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[5]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[31]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[4]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[4]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[30]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[3]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[3]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[29]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_negative_b[2]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_b[2]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  INVX0 U96 ( .INP(product_shift[28]), .ZN(n46) );
  INVX0 U97 ( .INP(n46), .ZN(n47) );
  NBUFFX2 U98 ( .INP(n51), .Z(n60) );
  NBUFFX2 U99 ( .INP(n50), .Z(n61) );
  NBUFFX2 U100 ( .INP(n51), .Z(n62) );
  NBUFFX2 U101 ( .INP(n50), .Z(n63) );
  NBUFFX2 U102 ( .INP(n51), .Z(n64) );
  NBUFFX2 U103 ( .INP(n50), .Z(n65) );
  NBUFFX2 U104 ( .INP(n51), .Z(n66) );
  NBUFFX2 U105 ( .INP(n50), .Z(n67) );
  NBUFFX2 U106 ( .INP(n51), .Z(n68) );
  NBUFFX2 U107 ( .INP(n51), .Z(n69) );
  NBUFFX2 U108 ( .INP(n50), .Z(n70) );
  NBUFFX2 U109 ( .INP(n74), .Z(n58) );
  NBUFFX2 U110 ( .INP(n74), .Z(n57) );
  NBUFFX2 U111 ( .INP(n74), .Z(n56) );
  NBUFFX2 U112 ( .INP(n74), .Z(n59) );
  NBUFFX2 U113 ( .INP(n72), .Z(n52) );
  NBUFFX2 U114 ( .INP(n72), .Z(n53) );
  NBUFFX2 U115 ( .INP(n73), .Z(n55) );
  NBUFFX2 U116 ( .INP(n73), .Z(n54) );
  NBUFFX2 U117 ( .INP(reset), .Z(n51) );
  NBUFFX2 U118 ( .INP(reset), .Z(n50) );
  NOR2X0 U119 ( .IN1(n71), .IN2(product_shift[1]), .QN(n74) );
  INVX0 U120 ( .INP(product_shift[0]), .ZN(n71) );
  INVX0 U122 ( .INP(product_shift[27]), .ZN(n48) );
  INVX0 U123 ( .INP(n48), .ZN(n49) );
endmodule


module booth6_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n38), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  XOR3X1 U1 ( .IN1(carry[38]), .IN2(B[38]), .IN3(A[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(carry[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[38]), .IN2(A[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[39]) );
  NAND3X1 U6 ( .IN1(n26), .IN2(n25), .IN3(n24), .QN(n15) );
  NAND3X1 U7 ( .IN1(n29), .IN2(n30), .IN3(n28), .QN(n11) );
  XOR2X1 U8 ( .IN1(n34), .IN2(carry[47]), .Q(SUM[47]) );
  XOR3X1 U9 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X1 U10 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U11 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U12 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U13 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U14 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U15 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U16 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U17 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U18 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U19 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  XOR3X1 U20 ( .IN1(n11), .IN2(B[45]), .IN3(A[45]), .Q(SUM[45]) );
  NAND2X0 U21 ( .IN1(A[45]), .IN2(carry[45]), .QN(n12) );
  NAND2X0 U22 ( .IN1(B[45]), .IN2(carry[45]), .QN(n13) );
  NAND2X0 U23 ( .IN1(B[45]), .IN2(A[45]), .QN(n14) );
  NAND3X0 U24 ( .IN1(n12), .IN2(n14), .IN3(n13), .QN(carry[46]) );
  DELLN2X2 U25 ( .INP(carry[41]), .Z(n16) );
  XOR3X2 U26 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  XOR3X2 U27 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U28 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U29 ( .IN1(A[40]), .IN2(B[40]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[40]), .IN2(carry[40]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[40]), .IN2(carry[40]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n19), .IN2(n18), .IN3(n17), .QN(carry[41]) );
  XOR2X1 U33 ( .IN1(A[41]), .IN2(B[41]), .Q(n20) );
  XOR2X1 U34 ( .IN1(n20), .IN2(n16), .Q(SUM[41]) );
  NAND2X0 U35 ( .IN1(A[41]), .IN2(B[41]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[41]), .IN2(carry[41]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[41]), .IN2(carry[41]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[42]) );
  NAND2X0 U39 ( .IN1(A[43]), .IN2(B[43]), .QN(n24) );
  NAND2X0 U40 ( .IN1(A[43]), .IN2(carry[43]), .QN(n25) );
  NAND2X0 U41 ( .IN1(B[43]), .IN2(carry[43]), .QN(n26) );
  NAND3X0 U42 ( .IN1(n26), .IN2(n25), .IN3(n24), .QN(carry[44]) );
  XOR2X1 U43 ( .IN1(A[44]), .IN2(B[44]), .Q(n27) );
  XOR2X1 U44 ( .IN1(n27), .IN2(n15), .Q(SUM[44]) );
  NAND2X0 U45 ( .IN1(A[44]), .IN2(B[44]), .QN(n28) );
  NAND2X0 U46 ( .IN1(A[44]), .IN2(carry[44]), .QN(n29) );
  NAND2X0 U47 ( .IN1(B[44]), .IN2(carry[44]), .QN(n30) );
  NAND3X0 U48 ( .IN1(n29), .IN2(n30), .IN3(n28), .QN(carry[45]) );
  NAND2X0 U49 ( .IN1(A[46]), .IN2(B[46]), .QN(n31) );
  NAND2X0 U50 ( .IN1(A[46]), .IN2(carry[46]), .QN(n32) );
  NAND2X0 U51 ( .IN1(B[46]), .IN2(carry[46]), .QN(n33) );
  NAND3X0 U52 ( .IN1(n33), .IN2(n32), .IN3(n31), .QN(carry[47]) );
  XOR2X1 U53 ( .IN1(A[47]), .IN2(B[47]), .Q(n34) );
  NAND2X0 U54 ( .IN1(A[47]), .IN2(B[47]), .QN(n35) );
  NAND2X0 U55 ( .IN1(A[47]), .IN2(carry[47]), .QN(n36) );
  NAND2X0 U56 ( .IN1(B[47]), .IN2(carry[47]), .QN(n37) );
  NAND3X0 U57 ( .IN1(n36), .IN2(n37), .IN3(n35), .QN(carry[48]) );
  AND2X1 U58 ( .IN1(A[26]), .IN2(B[26]), .Q(n38) );
  XOR2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_18_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n8), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n25), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR3X1 U6 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U7 ( .IN1(A[46]), .IN2(carry[46]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[46]), .IN2(carry[46]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[46]), .IN2(A[46]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[47]) );
  INVX0 U11 ( .INP(A[34]), .ZN(n7) );
  INVX0 U12 ( .INP(n7), .ZN(n8) );
  DELLN1X2 U13 ( .INP(carry[48]), .Z(n9) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n10) );
  XNOR2X1 U15 ( .IN1(n11), .IN2(n10), .Q(SUM[45]) );
  XNOR2X1 U16 ( .IN1(A[45]), .IN2(B[45]), .Q(n11) );
  XNOR2X1 U17 ( .IN1(n12), .IN2(n9), .Q(SUM[48]) );
  XNOR2X1 U18 ( .IN1(A[48]), .IN2(B[48]), .Q(n12) );
  XOR3X2 U19 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(B[44]), .QN(n13) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(carry[44]), .QN(n14) );
  NAND2X0 U22 ( .IN1(B[44]), .IN2(carry[44]), .QN(n15) );
  NAND3X0 U23 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[45]) );
  NAND2X0 U24 ( .IN1(A[45]), .IN2(B[45]), .QN(n16) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(carry[45]), .QN(n17) );
  NAND2X0 U26 ( .IN1(B[45]), .IN2(carry[45]), .QN(n18) );
  NAND3X0 U27 ( .IN1(n17), .IN2(n18), .IN3(n16), .QN(carry[46]) );
  XOR3X2 U28 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U32 ( .IN1(n21), .IN2(n20), .IN3(n19), .QN(carry[48]) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(B[48]), .QN(n22) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(carry[48]), .QN(n23) );
  NAND2X0 U35 ( .IN1(B[48]), .IN2(carry[48]), .QN(n24) );
  NAND3X0 U36 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[49]) );
  AND2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  XOR2X1 U38 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_18 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[18] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n73), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n73), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n51), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n50), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n45), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n43), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n65), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n63), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n63), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n63), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n63), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n63), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n63), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n63), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n63), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n63), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n63), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n58), .IN3(N75), .IN4(n54), .IN5(
        product_shift[9]), .IN6(n52), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n58), .IN3(N74), .IN4(n54), .IN5(
        product_shift[8]), .IN6(n53), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n58), .IN3(N73), .IN4(n54), .IN5(
        product_shift[7]), .IN6(n53), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n58), .IN3(N72), .IN4(n54), .IN5(
        product_shift[6]), .IN6(n53), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n58), .IN3(N71), .IN4(n54), .IN5(
        product_shift[5]), .IN6(n53), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n58), .IN3(N116), .IN4(n54), .IN5(
        product_shift[49]), .IN6(n53), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n58), .IN3(N70), .IN4(n54), .IN5(
        product_shift[4]), .IN6(n53), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n58), .IN3(N115), .IN4(n54), .IN5(
        product_shift[49]), .IN6(n53), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n58), .IN3(N114), .IN4(n54), .IN5(
        product_shift[48]), .IN6(n53), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n58), .IN3(N113), .IN4(n54), .IN5(
        product_shift[47]), .IN6(n53), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n58), .IN3(N112), .IN4(n54), .IN5(
        product_shift[46]), .IN6(n53), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n58), .IN3(N111), .IN4(n54), .IN5(
        product_shift[45]), .IN6(n53), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n59), .IN3(N110), .IN4(n55), .IN5(
        product_shift[44]), .IN6(n53), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n59), .IN3(N109), .IN4(n55), .IN5(
        product_shift[43]), .IN6(n75), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n59), .IN3(N108), .IN4(n55), .IN5(
        product_shift[42]), .IN6(n53), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n59), .IN3(N107), .IN4(n55), .IN5(
        product_shift[41]), .IN6(n52), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n59), .IN3(N106), .IN4(n55), .IN5(
        product_shift[40]), .IN6(n75), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n59), .IN3(N69), .IN4(n55), .IN5(
        product_shift[3]), .IN6(n75), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n59), .IN3(N105), .IN4(n55), .IN5(
        product_shift[39]), .IN6(n75), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n59), .IN3(N104), .IN4(n55), .IN5(
        product_shift[38]), .IN6(n75), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n59), .IN3(N103), .IN4(n55), .IN5(
        product_shift[37]), .IN6(n75), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n59), .IN3(N102), .IN4(n55), .IN5(
        product_shift[36]), .IN6(n75), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n59), .IN3(N101), .IN4(n55), .IN5(
        product_shift[35]), .IN6(n75), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n59), .IN3(N100), .IN4(n55), .IN5(
        product_shift[34]), .IN6(n75), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n60), .IN3(N99), .IN4(n55), .IN5(n11), .IN6(
        n53), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n60), .IN3(N98), .IN4(n57), .IN5(n17), .IN6(
        n75), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n60), .IN3(N97), .IN4(n56), .IN5(n23), .IN6(
        n75), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n60), .IN3(N96), .IN4(n57), .IN5(n29), .IN6(
        n75), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n60), .IN3(N68), .IN4(n57), .IN5(
        product_shift[2]), .IN6(n75), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n60), .IN3(N95), .IN4(n57), .IN5(n35), .IN6(
        n75), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n60), .IN3(N94), .IN4(n57), .IN5(n41), .IN6(
        n75), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n60), .IN3(N93), .IN4(n57), .IN5(n47), .IN6(
        n75), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n60), .IN3(N92), .IN4(n57), .IN5(n49), .IN6(
        n75), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n60), .IN3(N91), .IN4(n57), .IN5(
        product_shift[25]), .IN6(n75), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n60), .IN3(N90), .IN4(n57), .IN5(
        product_shift[24]), .IN6(n75), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n60), .IN3(N89), .IN4(n57), .IN5(
        product_shift[23]), .IN6(n52), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n61), .IN3(N88), .IN4(n56), .IN5(
        product_shift[22]), .IN6(n75), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n61), .IN3(N87), .IN4(n56), .IN5(
        product_shift[21]), .IN6(n52), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n61), .IN3(N86), .IN4(n56), .IN5(
        product_shift[20]), .IN6(n52), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n61), .IN3(N67), .IN4(n56), .IN5(n52), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n61), .IN3(N85), .IN4(n56), .IN5(
        product_shift[19]), .IN6(n52), .Q(product2[19]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n61), .IN3(N83), .IN4(n56), .IN5(
        product_shift[17]), .IN6(n52), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n61), .IN3(N82), .IN4(n56), .IN5(
        product_shift[16]), .IN6(n52), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n61), .IN3(N81), .IN4(n56), .IN5(
        product_shift[15]), .IN6(n52), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n61), .IN3(N80), .IN4(n56), .IN5(
        product_shift[14]), .IN6(n52), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n61), .IN3(N79), .IN4(n56), .IN5(
        product_shift[13]), .IN6(n52), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n61), .IN3(N78), .IN4(n56), .IN5(
        product_shift[12]), .IN6(n52), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n62), .IN3(N77), .IN4(n57), .IN5(
        product_shift[11]), .IN6(n52), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n62), .IN3(N76), .IN4(n57), .IN5(
        product_shift[10]), .IN6(n53), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n75) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n74), .Q(n76) );
  booth6_18_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, SYNOPSYS_UNCONNECTED__0, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_18_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, n45, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        SYNOPSYS_UNCONNECTED__2, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U48 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_negative_b[1]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_b[1]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  NBUFFX2 U96 ( .INP(n51), .Z(n63) );
  NBUFFX2 U97 ( .INP(n50), .Z(n64) );
  NBUFFX2 U98 ( .INP(n51), .Z(n65) );
  NBUFFX2 U99 ( .INP(n50), .Z(n66) );
  NBUFFX2 U100 ( .INP(n51), .Z(n67) );
  NBUFFX2 U101 ( .INP(n50), .Z(n68) );
  NBUFFX2 U102 ( .INP(n51), .Z(n69) );
  NBUFFX2 U103 ( .INP(n50), .Z(n70) );
  NBUFFX2 U104 ( .INP(n51), .Z(n71) );
  NBUFFX2 U105 ( .INP(n51), .Z(n72) );
  NBUFFX2 U106 ( .INP(n50), .Z(n73) );
  NBUFFX2 U107 ( .INP(n77), .Z(n60) );
  NBUFFX2 U108 ( .INP(n77), .Z(n59) );
  NBUFFX2 U109 ( .INP(n77), .Z(n58) );
  NBUFFX2 U110 ( .INP(n77), .Z(n61) );
  NBUFFX2 U111 ( .INP(n77), .Z(n62) );
  NBUFFX2 U112 ( .INP(n75), .Z(n52) );
  NBUFFX2 U113 ( .INP(n75), .Z(n53) );
  NBUFFX2 U114 ( .INP(n76), .Z(n55) );
  NBUFFX2 U115 ( .INP(n76), .Z(n54) );
  NBUFFX2 U116 ( .INP(n76), .Z(n56) );
  NBUFFX2 U117 ( .INP(n76), .Z(n57) );
  NBUFFX2 U118 ( .INP(reset), .Z(n51) );
  NBUFFX2 U119 ( .INP(reset), .Z(n50) );
  NOR2X0 U120 ( .IN1(n74), .IN2(product_shift[1]), .QN(n77) );
  INVX0 U121 ( .INP(product_shift[0]), .ZN(n74) );
  INVX0 U123 ( .INP(product_shift[27]), .ZN(n46) );
  INVX0 U124 ( .INP(n46), .ZN(n47) );
  INVX0 U125 ( .INP(product_shift[26]), .ZN(n48) );
  INVX0 U126 ( .INP(n48), .ZN(n49) );
endmodule


module booth6_17_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n40), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X2 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U6 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U8 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XOR3X1 U12 ( .IN1(A[48]), .IN2(B[48]), .IN3(n15), .Q(SUM[48]) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(B[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[48]), .IN2(carry[48]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[48]), .IN2(carry[48]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[49]) );
  XOR2X1 U17 ( .IN1(A[49]), .IN2(B[49]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(B[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[49]), .IN2(carry[49]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[49]), .IN2(carry[49]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[50]) );
  DELLN1X2 U23 ( .INP(carry[48]), .Z(n15) );
  DELLN2X2 U24 ( .INP(carry[44]), .Z(n16) );
  DELLN2X2 U25 ( .INP(carry[41]), .Z(n17) );
  DELLN2X2 U26 ( .INP(carry[47]), .Z(n18) );
  XOR3X2 U27 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  XOR3X2 U28 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U29 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U30 ( .IN1(A[40]), .IN2(B[40]), .QN(n19) );
  NAND2X0 U31 ( .IN1(A[40]), .IN2(carry[40]), .QN(n20) );
  NAND2X0 U32 ( .IN1(B[40]), .IN2(carry[40]), .QN(n21) );
  NAND3X0 U33 ( .IN1(n20), .IN2(n21), .IN3(n19), .QN(carry[41]) );
  XOR2X1 U34 ( .IN1(A[41]), .IN2(B[41]), .Q(n22) );
  XOR2X1 U35 ( .IN1(n22), .IN2(n17), .Q(SUM[41]) );
  NAND2X0 U36 ( .IN1(A[41]), .IN2(B[41]), .QN(n23) );
  NAND2X0 U37 ( .IN1(A[41]), .IN2(carry[41]), .QN(n24) );
  NAND2X0 U38 ( .IN1(B[41]), .IN2(carry[41]), .QN(n25) );
  NAND3X0 U39 ( .IN1(n24), .IN2(n25), .IN3(n23), .QN(carry[42]) );
  NAND2X0 U40 ( .IN1(A[43]), .IN2(B[43]), .QN(n26) );
  NAND2X0 U41 ( .IN1(A[43]), .IN2(carry[43]), .QN(n27) );
  NAND2X0 U42 ( .IN1(B[43]), .IN2(carry[43]), .QN(n28) );
  NAND3X0 U43 ( .IN1(n27), .IN2(n28), .IN3(n26), .QN(carry[44]) );
  XOR2X1 U44 ( .IN1(A[44]), .IN2(B[44]), .Q(n29) );
  XOR2X1 U45 ( .IN1(n29), .IN2(n16), .Q(SUM[44]) );
  NAND2X0 U46 ( .IN1(A[44]), .IN2(B[44]), .QN(n30) );
  NAND2X0 U47 ( .IN1(A[44]), .IN2(carry[44]), .QN(n31) );
  NAND2X0 U48 ( .IN1(B[44]), .IN2(carry[44]), .QN(n32) );
  NAND3X0 U49 ( .IN1(n31), .IN2(n32), .IN3(n30), .QN(carry[45]) );
  NAND2X0 U50 ( .IN1(A[46]), .IN2(B[46]), .QN(n33) );
  NAND2X0 U51 ( .IN1(A[46]), .IN2(carry[46]), .QN(n34) );
  NAND2X0 U52 ( .IN1(B[46]), .IN2(carry[46]), .QN(n35) );
  NAND3X0 U53 ( .IN1(n33), .IN2(n34), .IN3(n35), .QN(carry[47]) );
  XOR2X1 U54 ( .IN1(A[47]), .IN2(B[47]), .Q(n36) );
  XOR2X1 U55 ( .IN1(n36), .IN2(n18), .Q(SUM[47]) );
  NAND2X0 U56 ( .IN1(A[47]), .IN2(B[47]), .QN(n37) );
  NAND2X0 U57 ( .IN1(A[47]), .IN2(carry[47]), .QN(n38) );
  NAND2X0 U58 ( .IN1(B[47]), .IN2(carry[47]), .QN(n39) );
  NAND3X0 U59 ( .IN1(n38), .IN2(n39), .IN3(n37), .QN(carry[48]) );
  AND2X1 U60 ( .IN1(A[26]), .IN2(B[26]), .Q(n40) );
  XOR2X1 U61 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_17_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n8), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n25), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR3X1 U6 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U7 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  INVX0 U11 ( .INP(A[34]), .ZN(n7) );
  INVX0 U12 ( .INP(n7), .ZN(n8) );
  DELLN1X2 U13 ( .INP(carry[48]), .Z(n9) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n10) );
  XNOR2X1 U15 ( .IN1(n11), .IN2(n10), .Q(SUM[45]) );
  XNOR2X1 U16 ( .IN1(A[45]), .IN2(B[45]), .Q(n11) );
  XNOR2X1 U17 ( .IN1(n12), .IN2(n9), .Q(SUM[48]) );
  XNOR2X1 U18 ( .IN1(A[48]), .IN2(B[48]), .Q(n12) );
  XOR3X2 U19 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(B[44]), .QN(n13) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(carry[44]), .QN(n14) );
  NAND2X0 U22 ( .IN1(B[44]), .IN2(carry[44]), .QN(n15) );
  NAND3X0 U23 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[45]) );
  NAND2X0 U24 ( .IN1(A[45]), .IN2(B[45]), .QN(n16) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(carry[45]), .QN(n17) );
  NAND2X0 U26 ( .IN1(B[45]), .IN2(carry[45]), .QN(n18) );
  NAND3X0 U27 ( .IN1(n18), .IN2(n17), .IN3(n16), .QN(carry[46]) );
  XOR3X2 U28 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U32 ( .IN1(n20), .IN2(n21), .IN3(n19), .QN(carry[48]) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(B[48]), .QN(n22) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(carry[48]), .QN(n23) );
  NAND2X0 U35 ( .IN1(B[48]), .IN2(carry[48]), .QN(n24) );
  NAND3X0 U36 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[49]) );
  AND2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  XOR2X1 U38 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_17 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[17] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n70), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n70), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n45), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n43), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n62), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n61), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n59), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n59), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n59), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n59), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n59), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n59), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n59), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n59), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n59), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n59), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n55), .IN3(N75), .IN4(n53), .IN5(
        product_shift[9]), .IN6(n51), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n55), .IN3(N74), .IN4(n73), .IN5(
        product_shift[8]), .IN6(n52), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n55), .IN3(N73), .IN4(n73), .IN5(
        product_shift[7]), .IN6(n52), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n55), .IN3(N72), .IN4(n73), .IN5(
        product_shift[6]), .IN6(n52), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n55), .IN3(N71), .IN4(n73), .IN5(
        product_shift[5]), .IN6(n52), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n55), .IN3(N116), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n52), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n55), .IN3(N70), .IN4(n73), .IN5(
        product_shift[4]), .IN6(n52), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n55), .IN3(N115), .IN4(n73), .IN5(
        product_shift[49]), .IN6(n52), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n55), .IN3(N114), .IN4(n73), .IN5(
        product_shift[48]), .IN6(n52), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n55), .IN3(N113), .IN4(n73), .IN5(
        product_shift[47]), .IN6(n52), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n55), .IN3(N112), .IN4(n73), .IN5(
        product_shift[46]), .IN6(n52), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n55), .IN3(N111), .IN4(n73), .IN5(
        product_shift[45]), .IN6(n52), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n56), .IN3(N110), .IN4(n73), .IN5(
        product_shift[44]), .IN6(n72), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n58), .IN3(N109), .IN4(n73), .IN5(
        product_shift[43]), .IN6(n72), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n57), .IN3(N108), .IN4(n73), .IN5(
        product_shift[42]), .IN6(n72), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n58), .IN3(N107), .IN4(n73), .IN5(
        product_shift[41]), .IN6(n72), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n58), .IN3(N106), .IN4(n73), .IN5(
        product_shift[40]), .IN6(n72), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n58), .IN3(N69), .IN4(n73), .IN5(
        product_shift[3]), .IN6(n72), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n58), .IN3(N105), .IN4(n73), .IN5(
        product_shift[39]), .IN6(n72), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n58), .IN3(N104), .IN4(n54), .IN5(
        product_shift[38]), .IN6(n51), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n58), .IN3(N103), .IN4(n53), .IN5(
        product_shift[37]), .IN6(n52), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n58), .IN3(N102), .IN4(n54), .IN5(
        product_shift[36]), .IN6(n51), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n58), .IN3(N101), .IN4(n53), .IN5(
        product_shift[35]), .IN6(n52), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n58), .IN3(N100), .IN4(n54), .IN5(
        product_shift[34]), .IN6(n52), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n56), .IN3(N99), .IN4(n73), .IN5(n11), .IN6(
        n72), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n56), .IN3(N98), .IN4(n54), .IN5(n17), .IN6(
        n72), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n56), .IN3(N97), .IN4(n53), .IN5(n23), .IN6(
        n72), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n56), .IN3(N96), .IN4(n54), .IN5(n29), .IN6(
        n72), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n56), .IN3(N68), .IN4(n54), .IN5(
        product_shift[2]), .IN6(n72), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n56), .IN3(N95), .IN4(n54), .IN5(n35), .IN6(
        n72), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n56), .IN3(N94), .IN4(n54), .IN5(n41), .IN6(
        n72), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n56), .IN3(N93), .IN4(n54), .IN5(n47), .IN6(
        n72), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n56), .IN3(N92), .IN4(n54), .IN5(n49), .IN6(
        n72), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n56), .IN3(N91), .IN4(n54), .IN5(
        product_shift[25]), .IN6(n72), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n56), .IN3(N90), .IN4(n54), .IN5(
        product_shift[24]), .IN6(n72), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n56), .IN3(N89), .IN4(n54), .IN5(
        product_shift[23]), .IN6(n72), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n57), .IN3(N88), .IN4(n53), .IN5(
        product_shift[22]), .IN6(n72), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n57), .IN3(N87), .IN4(n53), .IN5(
        product_shift[21]), .IN6(n51), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n57), .IN3(N86), .IN4(n53), .IN5(
        product_shift[20]), .IN6(n51), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n57), .IN3(N67), .IN4(n53), .IN5(n51), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n57), .IN3(N85), .IN4(n53), .IN5(
        product_shift[19]), .IN6(n51), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n57), .IN3(N84), .IN4(n53), .IN5(
        product_shift[18]), .IN6(n51), .Q(product2[18]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n57), .IN3(N82), .IN4(n53), .IN5(
        product_shift[16]), .IN6(n51), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n57), .IN3(N81), .IN4(n53), .IN5(
        product_shift[15]), .IN6(n51), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n57), .IN3(N80), .IN4(n53), .IN5(
        product_shift[14]), .IN6(n51), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n57), .IN3(N79), .IN4(n53), .IN5(
        product_shift[13]), .IN6(n51), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n57), .IN3(N78), .IN4(n53), .IN5(
        product_shift[12]), .IN6(n51), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n58), .IN3(N77), .IN4(n54), .IN5(
        product_shift[11]), .IN6(n51), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n58), .IN3(N76), .IN4(n54), .IN5(
        product_shift[10]), .IN6(n52), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n72) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n71), .Q(n73) );
  booth6_17_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, SYNOPSYS_UNCONNECTED__0, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_17_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, n45, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        SYNOPSYS_UNCONNECTED__2, N31, N30, N29, N28, N27, N26, N25, N24, N23, 
        N22, N21, N20, N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U49 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_negative_b[1]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_b[1]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  NBUFFX2 U96 ( .INP(n50), .Z(n59) );
  NBUFFX2 U97 ( .INP(n50), .Z(n60) );
  NBUFFX2 U98 ( .INP(n50), .Z(n61) );
  NBUFFX2 U99 ( .INP(n50), .Z(n62) );
  NBUFFX2 U100 ( .INP(n50), .Z(n63) );
  NBUFFX2 U101 ( .INP(n50), .Z(n64) );
  NBUFFX2 U102 ( .INP(n50), .Z(n65) );
  NBUFFX2 U103 ( .INP(n50), .Z(n66) );
  NBUFFX2 U104 ( .INP(n68), .Z(n67) );
  NBUFFX2 U105 ( .INP(n68), .Z(n69) );
  NBUFFX2 U106 ( .INP(n50), .Z(n70) );
  NBUFFX2 U107 ( .INP(n50), .Z(n68) );
  NBUFFX2 U108 ( .INP(n74), .Z(n56) );
  NBUFFX2 U109 ( .INP(n74), .Z(n55) );
  NBUFFX2 U110 ( .INP(n74), .Z(n57) );
  NBUFFX2 U111 ( .INP(n74), .Z(n58) );
  NBUFFX2 U112 ( .INP(n72), .Z(n51) );
  NBUFFX2 U113 ( .INP(n72), .Z(n52) );
  NBUFFX2 U114 ( .INP(n73), .Z(n53) );
  NBUFFX2 U115 ( .INP(n73), .Z(n54) );
  NBUFFX2 U116 ( .INP(reset), .Z(n50) );
  NOR2X0 U117 ( .IN1(n71), .IN2(product_shift[1]), .QN(n74) );
  INVX0 U118 ( .INP(product_shift[0]), .ZN(n71) );
  INVX0 U120 ( .INP(product_shift[27]), .ZN(n46) );
  INVX0 U121 ( .INP(n46), .ZN(n47) );
  INVX0 U122 ( .INP(product_shift[26]), .ZN(n48) );
  INVX0 U123 ( .INP(n48), .ZN(n49) );
endmodule


module booth6_16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n39), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X2 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U6 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U8 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XOR3X2 U12 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(B[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[48]), .IN2(carry[48]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[48]), .IN2(carry[48]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[49]) );
  XOR2X1 U17 ( .IN1(A[49]), .IN2(B[49]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(B[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[49]), .IN2(carry[49]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[49]), .IN2(carry[49]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[50]) );
  DELLN2X2 U23 ( .INP(carry[41]), .Z(n15) );
  DELLN2X2 U24 ( .INP(carry[44]), .Z(n16) );
  DELLN2X2 U25 ( .INP(carry[47]), .Z(n17) );
  XOR3X2 U26 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  XOR3X2 U27 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U28 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U29 ( .IN1(A[40]), .IN2(B[40]), .QN(n18) );
  NAND2X0 U30 ( .IN1(A[40]), .IN2(carry[40]), .QN(n19) );
  NAND2X0 U31 ( .IN1(B[40]), .IN2(carry[40]), .QN(n20) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[41]) );
  XOR2X1 U33 ( .IN1(A[41]), .IN2(B[41]), .Q(n21) );
  XOR2X1 U34 ( .IN1(n21), .IN2(n15), .Q(SUM[41]) );
  NAND2X0 U35 ( .IN1(A[41]), .IN2(B[41]), .QN(n22) );
  NAND2X0 U36 ( .IN1(A[41]), .IN2(carry[41]), .QN(n23) );
  NAND2X0 U37 ( .IN1(B[41]), .IN2(carry[41]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[42]) );
  NAND2X0 U39 ( .IN1(A[43]), .IN2(B[43]), .QN(n25) );
  NAND2X0 U40 ( .IN1(A[43]), .IN2(carry[43]), .QN(n26) );
  NAND2X0 U41 ( .IN1(B[43]), .IN2(carry[43]), .QN(n27) );
  NAND3X0 U42 ( .IN1(n25), .IN2(n26), .IN3(n27), .QN(carry[44]) );
  XOR2X1 U43 ( .IN1(A[44]), .IN2(B[44]), .Q(n28) );
  XOR2X1 U44 ( .IN1(n28), .IN2(n16), .Q(SUM[44]) );
  NAND2X0 U45 ( .IN1(A[44]), .IN2(B[44]), .QN(n29) );
  NAND2X0 U46 ( .IN1(A[44]), .IN2(carry[44]), .QN(n30) );
  NAND2X0 U47 ( .IN1(B[44]), .IN2(carry[44]), .QN(n31) );
  NAND3X0 U48 ( .IN1(n31), .IN2(n30), .IN3(n29), .QN(carry[45]) );
  NAND2X0 U49 ( .IN1(A[46]), .IN2(B[46]), .QN(n32) );
  NAND2X0 U50 ( .IN1(A[46]), .IN2(carry[46]), .QN(n33) );
  NAND2X0 U51 ( .IN1(B[46]), .IN2(carry[46]), .QN(n34) );
  NAND3X0 U52 ( .IN1(n32), .IN2(n33), .IN3(n34), .QN(carry[47]) );
  XOR2X1 U53 ( .IN1(A[47]), .IN2(B[47]), .Q(n35) );
  XOR2X1 U54 ( .IN1(n35), .IN2(n17), .Q(SUM[47]) );
  NAND2X0 U55 ( .IN1(A[47]), .IN2(B[47]), .QN(n36) );
  NAND2X0 U56 ( .IN1(A[47]), .IN2(carry[47]), .QN(n37) );
  NAND2X0 U57 ( .IN1(B[47]), .IN2(carry[47]), .QN(n38) );
  NAND3X0 U58 ( .IN1(n38), .IN2(n37), .IN3(n36), .QN(carry[48]) );
  AND2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(n39) );
  XOR2X1 U60 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_16_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n26), .CO(carry[28]), .S(SUM[27])
         );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX2 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX2 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX2 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XNOR3X1 U1 ( .IN1(A[50]), .IN2(B[50]), .IN3(n1), .Q(SUM[50]) );
  AND3X1 U2 ( .IN1(n5), .IN2(n6), .IN3(n7), .Q(n1) );
  XOR3X1 U3 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U4 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X1 U5 ( .IN1(carry[37]), .IN2(B[37]), .IN3(A[37]), .Q(SUM[37]) );
  NAND2X1 U6 ( .IN1(A[37]), .IN2(carry[37]), .QN(n2) );
  NAND2X1 U7 ( .IN1(B[37]), .IN2(carry[37]), .QN(n3) );
  NAND2X1 U8 ( .IN1(B[37]), .IN2(A[37]), .QN(n4) );
  NAND3X0 U9 ( .IN1(n2), .IN2(n4), .IN3(n3), .QN(carry[38]) );
  XOR3X1 U10 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U11 ( .IN1(A[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U12 ( .IN1(B[49]), .IN2(carry[49]), .QN(n6) );
  NAND2X1 U13 ( .IN1(B[49]), .IN2(A[49]), .QN(n7) );
  INVX0 U14 ( .INP(A[34]), .ZN(n8) );
  INVX0 U15 ( .INP(n8), .ZN(n9) );
  DELLN1X2 U16 ( .INP(carry[48]), .Z(n10) );
  DELLN2X2 U17 ( .INP(carry[45]), .Z(n11) );
  XNOR2X1 U18 ( .IN1(n12), .IN2(n11), .Q(SUM[45]) );
  XNOR2X1 U19 ( .IN1(A[45]), .IN2(B[45]), .Q(n12) );
  XNOR2X1 U20 ( .IN1(n13), .IN2(n10), .Q(SUM[48]) );
  XNOR2X1 U21 ( .IN1(A[48]), .IN2(B[48]), .Q(n13) );
  NAND2X0 U22 ( .IN1(A[44]), .IN2(B[44]), .QN(n14) );
  NAND2X0 U23 ( .IN1(A[44]), .IN2(carry[44]), .QN(n15) );
  NAND2X0 U24 ( .IN1(B[44]), .IN2(carry[44]), .QN(n16) );
  NAND3X0 U25 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[45]) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(B[45]), .QN(n17) );
  NAND2X0 U27 ( .IN1(A[45]), .IN2(carry[45]), .QN(n18) );
  NAND2X0 U28 ( .IN1(B[45]), .IN2(carry[45]), .QN(n19) );
  NAND3X0 U29 ( .IN1(n18), .IN2(n19), .IN3(n17), .QN(carry[46]) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(B[47]), .QN(n20) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(carry[47]), .QN(n21) );
  NAND2X0 U32 ( .IN1(B[47]), .IN2(carry[47]), .QN(n22) );
  NAND3X0 U33 ( .IN1(n21), .IN2(n22), .IN3(n20), .QN(carry[48]) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(B[48]), .QN(n23) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(carry[48]), .QN(n24) );
  NAND2X0 U36 ( .IN1(B[48]), .IN2(carry[48]), .QN(n25) );
  NAND3X0 U37 ( .IN1(n24), .IN2(n25), .IN3(n23), .QN(carry[49]) );
  AND2X1 U38 ( .IN1(A[26]), .IN2(B[26]), .Q(n26) );
  XOR2X1 U39 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_16 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[16] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n76), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n76), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n45), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n69), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n69), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n69), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n69), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n43), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n68), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n67), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n65), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n65), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n65), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n65), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n65), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n65), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n65), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n65), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n65), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n65), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n60), .IN3(N75), .IN4(n55), .IN5(
        product_shift[9]), .IN6(n51), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n60), .IN3(N74), .IN4(n55), .IN5(
        product_shift[8]), .IN6(n54), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n60), .IN3(N73), .IN4(n55), .IN5(
        product_shift[7]), .IN6(n54), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n60), .IN3(N72), .IN4(n55), .IN5(
        product_shift[6]), .IN6(n54), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n60), .IN3(N71), .IN4(n55), .IN5(
        product_shift[5]), .IN6(n54), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(n60), .IN2(N65), .IN3(N116), .IN4(n55), .IN5(
        product_shift[49]), .IN6(n54), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n60), .IN3(N70), .IN4(n55), .IN5(
        product_shift[4]), .IN6(n54), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n60), .IN3(N115), .IN4(n55), .IN5(
        product_shift[49]), .IN6(n54), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n60), .IN3(N114), .IN4(n55), .IN5(
        product_shift[48]), .IN6(n54), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n60), .IN3(N113), .IN4(n55), .IN5(
        product_shift[47]), .IN6(n54), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n60), .IN3(N112), .IN4(n55), .IN5(
        product_shift[46]), .IN6(n54), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n60), .IN3(N111), .IN4(n55), .IN5(
        product_shift[45]), .IN6(n54), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n61), .IN3(N110), .IN4(n56), .IN5(
        product_shift[44]), .IN6(n53), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n61), .IN3(N109), .IN4(n56), .IN5(
        product_shift[43]), .IN6(n53), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n61), .IN3(N108), .IN4(n56), .IN5(
        product_shift[42]), .IN6(n53), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n61), .IN3(N107), .IN4(n56), .IN5(
        product_shift[41]), .IN6(n53), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n61), .IN3(N106), .IN4(n56), .IN5(
        product_shift[40]), .IN6(n53), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n61), .IN3(N69), .IN4(n56), .IN5(
        product_shift[3]), .IN6(n53), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n61), .IN3(N105), .IN4(n56), .IN5(
        product_shift[39]), .IN6(n53), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n61), .IN3(N104), .IN4(n56), .IN5(
        product_shift[38]), .IN6(n53), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n61), .IN3(N103), .IN4(n56), .IN5(
        product_shift[37]), .IN6(n53), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n61), .IN3(N102), .IN4(n56), .IN5(
        product_shift[36]), .IN6(n53), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n61), .IN3(N101), .IN4(n56), .IN5(
        product_shift[35]), .IN6(n53), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n61), .IN3(N100), .IN4(n56), .IN5(
        product_shift[34]), .IN6(n53), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n62), .IN3(N99), .IN4(n57), .IN5(n11), .IN6(
        n53), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n62), .IN3(N98), .IN4(n57), .IN5(n17), .IN6(
        n52), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n62), .IN3(N97), .IN4(n57), .IN5(n23), .IN6(
        n52), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n62), .IN3(N96), .IN4(n57), .IN5(n29), .IN6(
        n52), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n62), .IN3(N68), .IN4(n57), .IN5(
        product_shift[2]), .IN6(n52), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n62), .IN3(N95), .IN4(n57), .IN5(n35), .IN6(
        n52), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n62), .IN3(N94), .IN4(n57), .IN5(n41), .IN6(
        n52), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n62), .IN3(N93), .IN4(n57), .IN5(n47), .IN6(
        n52), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n62), .IN3(N92), .IN4(n57), .IN5(n49), .IN6(
        n52), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n62), .IN3(N91), .IN4(n57), .IN5(
        product_shift[25]), .IN6(n52), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n62), .IN3(N90), .IN4(n57), .IN5(
        product_shift[24]), .IN6(n52), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n62), .IN3(N89), .IN4(n57), .IN5(
        product_shift[23]), .IN6(n52), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n63), .IN3(N88), .IN4(n58), .IN5(
        product_shift[22]), .IN6(n52), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n63), .IN3(N87), .IN4(n58), .IN5(
        product_shift[21]), .IN6(n51), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n63), .IN3(N86), .IN4(n58), .IN5(
        product_shift[20]), .IN6(n51), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n63), .IN3(N67), .IN4(n58), .IN5(n51), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n63), .IN3(N85), .IN4(n58), .IN5(
        product_shift[19]), .IN6(n51), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n63), .IN3(N84), .IN4(n58), .IN5(
        product_shift[18]), .IN6(n51), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n63), .IN3(N83), .IN4(n58), .IN5(
        product_shift[17]), .IN6(n51), .Q(product2[17]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n63), .IN3(N81), .IN4(n58), .IN5(
        product_shift[15]), .IN6(n51), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n63), .IN3(N80), .IN4(n58), .IN5(
        product_shift[14]), .IN6(n51), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n63), .IN3(N79), .IN4(n58), .IN5(
        product_shift[13]), .IN6(n51), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n63), .IN3(N78), .IN4(n58), .IN5(
        product_shift[12]), .IN6(n51), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n64), .IN3(N77), .IN4(n59), .IN5(
        product_shift[11]), .IN6(n51), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n64), .IN3(N76), .IN4(n59), .IN5(
        product_shift[10]), .IN6(n52), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n78) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n77), .Q(n79) );
  booth6_16_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, SYNOPSYS_UNCONNECTED__0, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_16_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, n45, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        SYNOPSYS_UNCONNECTED__2, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U50 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_negative_b[1]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_b[1]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  NBUFFX2 U96 ( .INP(n50), .Z(n65) );
  NBUFFX2 U97 ( .INP(n50), .Z(n66) );
  NBUFFX2 U98 ( .INP(n50), .Z(n67) );
  NBUFFX2 U99 ( .INP(n50), .Z(n68) );
  NBUFFX2 U100 ( .INP(n50), .Z(n69) );
  NBUFFX2 U101 ( .INP(n50), .Z(n70) );
  NBUFFX2 U102 ( .INP(n50), .Z(n71) );
  NBUFFX2 U103 ( .INP(n50), .Z(n72) );
  NBUFFX2 U104 ( .INP(n50), .Z(n74) );
  NBUFFX2 U105 ( .INP(n50), .Z(n75) );
  NBUFFX2 U106 ( .INP(n50), .Z(n76) );
  NBUFFX2 U107 ( .INP(n50), .Z(n73) );
  NBUFFX2 U108 ( .INP(n80), .Z(n62) );
  NBUFFX2 U109 ( .INP(n80), .Z(n61) );
  NBUFFX2 U110 ( .INP(n80), .Z(n60) );
  NBUFFX2 U111 ( .INP(n80), .Z(n63) );
  NBUFFX2 U112 ( .INP(n80), .Z(n64) );
  NBUFFX2 U113 ( .INP(n78), .Z(n52) );
  NBUFFX2 U114 ( .INP(n78), .Z(n53) );
  NBUFFX2 U115 ( .INP(n78), .Z(n51) );
  NBUFFX2 U116 ( .INP(n78), .Z(n54) );
  NBUFFX2 U117 ( .INP(n79), .Z(n57) );
  NBUFFX2 U118 ( .INP(n79), .Z(n56) );
  NBUFFX2 U119 ( .INP(n79), .Z(n55) );
  NBUFFX2 U120 ( .INP(n79), .Z(n58) );
  NBUFFX2 U121 ( .INP(n79), .Z(n59) );
  NBUFFX2 U122 ( .INP(reset), .Z(n50) );
  NOR2X0 U123 ( .IN1(n77), .IN2(product_shift[1]), .QN(n80) );
  INVX0 U124 ( .INP(product_shift[0]), .ZN(n77) );
  INVX0 U126 ( .INP(product_shift[27]), .ZN(n46) );
  INVX0 U127 ( .INP(n46), .ZN(n47) );
  INVX0 U128 ( .INP(product_shift[26]), .ZN(n48) );
  INVX0 U129 ( .INP(n48), .ZN(n49) );
endmodule


module booth6_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X2 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U6 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U8 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XOR3X2 U12 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(B[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[48]), .IN2(carry[48]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[48]), .IN2(carry[48]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[49]) );
  XOR2X1 U17 ( .IN1(A[49]), .IN2(B[49]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(B[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[49]), .IN2(carry[49]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[49]), .IN2(carry[49]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[50]) );
  DELLN2X2 U23 ( .INP(carry[41]), .Z(n15) );
  DELLN2X2 U24 ( .INP(carry[47]), .Z(n16) );
  DELLN2X2 U25 ( .INP(carry[44]), .Z(n17) );
  AND2X1 U26 ( .IN1(A[26]), .IN2(B[26]), .Q(n42) );
  XOR3X1 U27 ( .IN1(B[27]), .IN2(n42), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U28 ( .IN1(n42), .IN2(B[27]), .QN(n40) );
  XOR3X1 U29 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X1 U30 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  XOR3X1 U31 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U32 ( .IN1(A[40]), .IN2(B[40]), .QN(n18) );
  NAND2X0 U33 ( .IN1(A[40]), .IN2(carry[40]), .QN(n19) );
  NAND2X0 U34 ( .IN1(B[40]), .IN2(carry[40]), .QN(n20) );
  NAND3X0 U35 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[41]) );
  XOR2X1 U36 ( .IN1(A[41]), .IN2(B[41]), .Q(n21) );
  XOR2X1 U37 ( .IN1(n21), .IN2(n15), .Q(SUM[41]) );
  NAND2X0 U38 ( .IN1(A[41]), .IN2(B[41]), .QN(n22) );
  NAND2X0 U39 ( .IN1(A[41]), .IN2(carry[41]), .QN(n23) );
  NAND2X0 U40 ( .IN1(B[41]), .IN2(carry[41]), .QN(n24) );
  NAND3X0 U41 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[42]) );
  NAND2X0 U42 ( .IN1(A[43]), .IN2(B[43]), .QN(n25) );
  NAND2X0 U43 ( .IN1(A[43]), .IN2(carry[43]), .QN(n26) );
  NAND2X0 U44 ( .IN1(B[43]), .IN2(carry[43]), .QN(n27) );
  NAND3X0 U45 ( .IN1(n25), .IN2(n26), .IN3(n27), .QN(carry[44]) );
  XOR2X1 U46 ( .IN1(A[44]), .IN2(B[44]), .Q(n28) );
  XOR2X1 U47 ( .IN1(n28), .IN2(n17), .Q(SUM[44]) );
  NAND2X0 U48 ( .IN1(A[44]), .IN2(B[44]), .QN(n29) );
  NAND2X0 U49 ( .IN1(A[44]), .IN2(carry[44]), .QN(n30) );
  NAND2X0 U50 ( .IN1(B[44]), .IN2(carry[44]), .QN(n31) );
  NAND3X0 U51 ( .IN1(n31), .IN2(n30), .IN3(n29), .QN(carry[45]) );
  NAND2X0 U52 ( .IN1(A[46]), .IN2(B[46]), .QN(n32) );
  NAND2X0 U53 ( .IN1(A[46]), .IN2(carry[46]), .QN(n33) );
  NAND2X0 U54 ( .IN1(B[46]), .IN2(carry[46]), .QN(n34) );
  NAND3X0 U55 ( .IN1(n32), .IN2(n33), .IN3(n34), .QN(carry[47]) );
  XOR2X1 U56 ( .IN1(A[47]), .IN2(B[47]), .Q(n35) );
  XOR2X1 U57 ( .IN1(n35), .IN2(n16), .Q(SUM[47]) );
  NAND2X0 U58 ( .IN1(A[47]), .IN2(B[47]), .QN(n36) );
  NAND2X0 U59 ( .IN1(A[47]), .IN2(carry[47]), .QN(n37) );
  NAND2X0 U60 ( .IN1(B[47]), .IN2(carry[47]), .QN(n38) );
  NAND3X0 U61 ( .IN1(n37), .IN2(n38), .IN3(n36), .QN(carry[48]) );
  NAND2X0 U62 ( .IN1(A[27]), .IN2(B[27]), .QN(n39) );
  NAND2X0 U63 ( .IN1(n42), .IN2(A[27]), .QN(n41) );
  NAND3X0 U64 ( .IN1(n39), .IN2(n41), .IN3(n40), .QN(carry[28]) );
  XOR2X1 U65 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_15_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR2X1 U6 ( .IN1(n21), .IN2(n7), .Q(SUM[48]) );
  XOR3X1 U7 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U8 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  DELLN1X2 U12 ( .INP(carry[48]), .Z(n7) );
  XOR3X1 U13 ( .IN1(B[27]), .IN2(n28), .IN3(A[27]), .Q(SUM[27]) );
  INVX0 U14 ( .INP(A[34]), .ZN(n8) );
  INVX0 U15 ( .INP(n8), .ZN(n9) );
  DELLN2X2 U16 ( .INP(carry[45]), .Z(n10) );
  NAND2X0 U17 ( .IN1(n28), .IN2(B[27]), .QN(n26) );
  XOR3X2 U18 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n11) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n12) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n13) );
  NAND3X0 U22 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n14) );
  XOR2X1 U24 ( .IN1(n14), .IN2(n10), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n16) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[46]) );
  XOR3X2 U29 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(B[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(carry[47]), .QN(n19) );
  NAND2X0 U32 ( .IN1(B[47]), .IN2(carry[47]), .QN(n20) );
  NAND3X0 U33 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[48]) );
  XOR2X1 U34 ( .IN1(A[48]), .IN2(B[48]), .Q(n21) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n22) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n23) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n23), .IN2(n24), .IN3(n22), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n25) );
  NAND2X0 U40 ( .IN1(n28), .IN2(A[27]), .QN(n27) );
  NAND3X0 U41 ( .IN1(n25), .IN2(n27), .IN3(n26), .QN(carry[28]) );
  AND2X4 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(n28) );
  XOR2X1 U43 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_15 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[15] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n64), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n64), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n60), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n60), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n60), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n60), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n59), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n58), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n58), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n58), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n58), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n58), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n57), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n57), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n57), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n56), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n56), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n56), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n56), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n56), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n56), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n55), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n55), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n55), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n55), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n53), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n53), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n53), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n53), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n53), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n53), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n53), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n53), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n53), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n53), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n53), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n53), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n49), .IN3(N75), .IN4(n47), .IN5(
        product_shift[9]), .IN6(n45), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n49), .IN3(N74), .IN4(n67), .IN5(
        product_shift[8]), .IN6(n46), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n49), .IN3(N73), .IN4(n67), .IN5(
        product_shift[7]), .IN6(n46), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n49), .IN3(N72), .IN4(n67), .IN5(
        product_shift[6]), .IN6(n46), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n49), .IN3(N71), .IN4(n67), .IN5(
        product_shift[5]), .IN6(n46), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n49), .IN3(N116), .IN4(n67), .IN5(
        product_shift[49]), .IN6(n46), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n49), .IN3(N70), .IN4(n67), .IN5(
        product_shift[4]), .IN6(n46), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n49), .IN3(N115), .IN4(n67), .IN5(
        product_shift[49]), .IN6(n46), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n49), .IN3(N114), .IN4(n67), .IN5(
        product_shift[48]), .IN6(n46), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n49), .IN3(N113), .IN4(n67), .IN5(
        product_shift[47]), .IN6(n46), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n49), .IN3(N112), .IN4(n67), .IN5(
        product_shift[46]), .IN6(n46), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n49), .IN3(N111), .IN4(n67), .IN5(
        product_shift[45]), .IN6(n46), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n50), .IN3(N110), .IN4(n67), .IN5(
        product_shift[44]), .IN6(n66), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n52), .IN3(N109), .IN4(n67), .IN5(
        product_shift[43]), .IN6(n66), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n51), .IN3(N108), .IN4(n67), .IN5(
        product_shift[42]), .IN6(n66), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n52), .IN3(N107), .IN4(n67), .IN5(
        product_shift[41]), .IN6(n66), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n52), .IN3(N106), .IN4(n67), .IN5(
        product_shift[40]), .IN6(n66), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n52), .IN3(N69), .IN4(n67), .IN5(
        product_shift[3]), .IN6(n66), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n52), .IN3(N105), .IN4(n67), .IN5(
        product_shift[39]), .IN6(n66), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n52), .IN3(N104), .IN4(n48), .IN5(
        product_shift[38]), .IN6(n45), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n52), .IN3(N103), .IN4(n47), .IN5(
        product_shift[37]), .IN6(n46), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n52), .IN3(N102), .IN4(n48), .IN5(
        product_shift[36]), .IN6(n45), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n52), .IN3(N101), .IN4(n47), .IN5(
        product_shift[35]), .IN6(n46), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n52), .IN3(N100), .IN4(n48), .IN5(
        product_shift[34]), .IN6(n46), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n50), .IN3(N99), .IN4(n67), .IN5(n11), .IN6(
        n66), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n50), .IN3(N98), .IN4(n48), .IN5(n17), .IN6(
        n66), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n50), .IN3(N97), .IN4(n47), .IN5(n23), .IN6(
        n66), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n50), .IN3(N96), .IN4(n48), .IN5(n29), .IN6(
        n66), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n50), .IN3(N68), .IN4(n48), .IN5(
        product_shift[2]), .IN6(n66), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n50), .IN3(N95), .IN4(n48), .IN5(n35), .IN6(
        n66), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n50), .IN3(N94), .IN4(n48), .IN5(n41), .IN6(
        n66), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n50), .IN3(N93), .IN4(n48), .IN5(n43), .IN6(
        n66), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n50), .IN3(N92), .IN4(n48), .IN5(
        product_shift[26]), .IN6(n66), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n50), .IN3(N91), .IN4(n48), .IN5(
        product_shift[25]), .IN6(n66), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n50), .IN3(N90), .IN4(n48), .IN5(
        product_shift[24]), .IN6(n66), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n50), .IN3(N89), .IN4(n48), .IN5(
        product_shift[23]), .IN6(n66), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n51), .IN3(N88), .IN4(n47), .IN5(
        product_shift[22]), .IN6(n66), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n51), .IN3(N87), .IN4(n47), .IN5(
        product_shift[21]), .IN6(n45), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n51), .IN3(N86), .IN4(n47), .IN5(
        product_shift[20]), .IN6(n45), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n51), .IN3(N67), .IN4(n47), .IN5(n45), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n51), .IN3(N85), .IN4(n47), .IN5(
        product_shift[19]), .IN6(n45), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n51), .IN3(N84), .IN4(n47), .IN5(
        product_shift[18]), .IN6(n45), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n51), .IN3(N83), .IN4(n47), .IN5(
        product_shift[17]), .IN6(n45), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n51), .IN3(N82), .IN4(n47), .IN5(
        product_shift[16]), .IN6(n45), .Q(product2[16]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n51), .IN3(N80), .IN4(n47), .IN5(
        product_shift[14]), .IN6(n45), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n51), .IN3(N79), .IN4(n47), .IN5(
        product_shift[13]), .IN6(n45), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n51), .IN3(N78), .IN4(n47), .IN5(
        product_shift[12]), .IN6(n45), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n52), .IN3(N77), .IN4(n48), .IN5(
        product_shift[11]), .IN6(n45), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n52), .IN3(N76), .IN4(n48), .IN5(
        product_shift[10]), .IN6(n46), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n66) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n65), .Q(n67) );
  booth6_15_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, product_shift[26:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, 
        combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, SYNOPSYS_UNCONNECTED__0, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_15_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, product_shift[26:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        SYNOPSYS_UNCONNECTED__2, N29, N28, N27, N26, N25, N24, N23, N22, N21, 
        N20, N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U51 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  NBUFFX2 U92 ( .INP(n44), .Z(n53) );
  NBUFFX2 U93 ( .INP(n44), .Z(n54) );
  NBUFFX2 U94 ( .INP(n44), .Z(n55) );
  NBUFFX2 U95 ( .INP(n44), .Z(n56) );
  NBUFFX2 U96 ( .INP(n44), .Z(n57) );
  NBUFFX2 U97 ( .INP(n44), .Z(n58) );
  NBUFFX2 U98 ( .INP(n44), .Z(n59) );
  NBUFFX2 U99 ( .INP(n44), .Z(n60) );
  NBUFFX2 U100 ( .INP(n44), .Z(n62) );
  NBUFFX2 U101 ( .INP(n44), .Z(n63) );
  NBUFFX2 U102 ( .INP(n44), .Z(n64) );
  NBUFFX2 U103 ( .INP(n44), .Z(n61) );
  NBUFFX2 U104 ( .INP(n68), .Z(n50) );
  NBUFFX2 U105 ( .INP(n68), .Z(n49) );
  NBUFFX2 U106 ( .INP(n68), .Z(n51) );
  NBUFFX2 U107 ( .INP(n68), .Z(n52) );
  NBUFFX2 U108 ( .INP(n66), .Z(n45) );
  NBUFFX2 U109 ( .INP(n66), .Z(n46) );
  NBUFFX2 U110 ( .INP(n67), .Z(n47) );
  NBUFFX2 U111 ( .INP(n67), .Z(n48) );
  NBUFFX2 U112 ( .INP(reset), .Z(n44) );
  NOR2X0 U113 ( .IN1(n65), .IN2(product_shift[1]), .QN(n68) );
  INVX0 U114 ( .INP(product_shift[0]), .ZN(n65) );
  INVX0 U116 ( .INP(product_shift[27]), .ZN(n42) );
  INVX0 U117 ( .INP(n42), .ZN(n43) );
endmodule


module booth6_14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[45]), .IN2(B[45]), .IN3(A[45]), .Q(SUM[45]) );
  NAND2X0 U2 ( .IN1(A[45]), .IN2(carry[45]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[45]), .IN2(carry[45]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[45]), .IN2(A[45]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[46]) );
  XOR3X2 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U7 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U11 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U13 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  DELLN2X2 U17 ( .INP(carry[41]), .Z(n11) );
  DELLN2X2 U18 ( .INP(carry[47]), .Z(n12) );
  DELLN2X2 U19 ( .INP(carry[44]), .Z(n13) );
  AND2X1 U20 ( .IN1(A[26]), .IN2(B[26]), .Q(n38) );
  XOR3X1 U21 ( .IN1(B[27]), .IN2(n38), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U22 ( .IN1(n38), .IN2(B[27]), .QN(n36) );
  XOR3X1 U23 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X1 U24 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  XOR3X1 U25 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U26 ( .IN1(A[40]), .IN2(B[40]), .QN(n14) );
  NAND2X0 U27 ( .IN1(A[40]), .IN2(carry[40]), .QN(n15) );
  NAND2X0 U28 ( .IN1(B[40]), .IN2(carry[40]), .QN(n16) );
  NAND3X0 U29 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(carry[41]) );
  XOR2X1 U30 ( .IN1(A[41]), .IN2(B[41]), .Q(n17) );
  XOR2X1 U31 ( .IN1(n17), .IN2(n11), .Q(SUM[41]) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(B[41]), .QN(n18) );
  NAND2X0 U33 ( .IN1(A[41]), .IN2(carry[41]), .QN(n19) );
  NAND2X0 U34 ( .IN1(B[41]), .IN2(carry[41]), .QN(n20) );
  NAND3X0 U35 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[42]) );
  NAND2X0 U36 ( .IN1(A[43]), .IN2(B[43]), .QN(n21) );
  NAND2X0 U37 ( .IN1(A[43]), .IN2(carry[43]), .QN(n22) );
  NAND2X0 U38 ( .IN1(B[43]), .IN2(carry[43]), .QN(n23) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n23), .IN3(n21), .QN(carry[44]) );
  XOR2X1 U40 ( .IN1(A[44]), .IN2(B[44]), .Q(n24) );
  XOR2X1 U41 ( .IN1(n24), .IN2(n13), .Q(SUM[44]) );
  NAND2X0 U42 ( .IN1(A[44]), .IN2(B[44]), .QN(n25) );
  NAND2X0 U43 ( .IN1(A[44]), .IN2(carry[44]), .QN(n26) );
  NAND2X0 U44 ( .IN1(B[44]), .IN2(carry[44]), .QN(n27) );
  NAND3X0 U45 ( .IN1(n26), .IN2(n27), .IN3(n25), .QN(carry[45]) );
  NAND2X0 U46 ( .IN1(A[46]), .IN2(B[46]), .QN(n28) );
  NAND2X0 U47 ( .IN1(A[46]), .IN2(carry[46]), .QN(n29) );
  NAND2X0 U48 ( .IN1(B[46]), .IN2(carry[46]), .QN(n30) );
  NAND3X0 U49 ( .IN1(n30), .IN2(n29), .IN3(n28), .QN(carry[47]) );
  XOR2X1 U50 ( .IN1(A[47]), .IN2(B[47]), .Q(n31) );
  XOR2X1 U51 ( .IN1(n31), .IN2(n12), .Q(SUM[47]) );
  NAND2X0 U52 ( .IN1(A[47]), .IN2(B[47]), .QN(n32) );
  NAND2X0 U53 ( .IN1(A[47]), .IN2(carry[47]), .QN(n33) );
  NAND2X0 U54 ( .IN1(B[47]), .IN2(carry[47]), .QN(n34) );
  NAND3X0 U55 ( .IN1(n33), .IN2(n34), .IN3(n32), .QN(carry[48]) );
  NAND2X0 U56 ( .IN1(A[27]), .IN2(B[27]), .QN(n35) );
  NAND2X0 U57 ( .IN1(n38), .IN2(A[27]), .QN(n37) );
  NAND3X0 U58 ( .IN1(n35), .IN2(n37), .IN3(n36), .QN(carry[28]) );
  XOR2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n8), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR2X1 U6 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  XOR3X1 U7 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U8 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  XOR3X1 U12 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  INVX0 U13 ( .INP(A[34]), .ZN(n7) );
  INVX0 U14 ( .INP(n7), .ZN(n8) );
  DELLN2X2 U15 ( .INP(carry[45]), .Z(n9) );
  NAND2X0 U16 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  XOR3X2 U17 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U18 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U20 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U21 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U22 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U23 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U24 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U26 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U27 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[46]) );
  XOR3X2 U28 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U36 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U37 ( .IN1(n23), .IN2(n22), .IN3(n21), .QN(carry[49]) );
  NAND2X0 U38 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U39 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U40 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  AND2X4 U41 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_14 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[14] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n65), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n65), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n61), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n60), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n16), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n22), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n28), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n34), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n40), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n59), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n58), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n58), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n58), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n5), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n14), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n20), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n26), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n32), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n38), .CLK(clk), .RSTB(n57), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n57), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n57), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n56), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n56), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n54), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n54), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n54), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n54), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n54), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n54), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n54), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n54), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n54), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n54), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n54), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n50), .IN3(N75), .IN4(n48), .IN5(
        product_shift[9]), .IN6(n46), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n50), .IN3(N74), .IN4(n68), .IN5(
        product_shift[8]), .IN6(n47), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n50), .IN3(N73), .IN4(n68), .IN5(
        product_shift[7]), .IN6(n47), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n50), .IN3(N72), .IN4(n68), .IN5(
        product_shift[6]), .IN6(n47), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n50), .IN3(N71), .IN4(n68), .IN5(
        product_shift[5]), .IN6(n47), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n50), .IN3(n68), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n47), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n50), .IN3(N70), .IN4(n68), .IN5(
        product_shift[4]), .IN6(n47), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n50), .IN3(N115), .IN4(n68), .IN5(
        product_shift[49]), .IN6(n47), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n50), .IN3(N114), .IN4(n68), .IN5(
        product_shift[48]), .IN6(n47), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n50), .IN3(N113), .IN4(n68), .IN5(
        product_shift[47]), .IN6(n47), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n50), .IN3(N112), .IN4(n68), .IN5(
        product_shift[46]), .IN6(n47), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n50), .IN3(N111), .IN4(n68), .IN5(
        product_shift[45]), .IN6(n47), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n51), .IN3(N110), .IN4(n68), .IN5(
        product_shift[44]), .IN6(n67), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n53), .IN3(N109), .IN4(n68), .IN5(
        product_shift[43]), .IN6(n67), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n52), .IN3(N108), .IN4(n68), .IN5(
        product_shift[42]), .IN6(n67), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n53), .IN3(N107), .IN4(n68), .IN5(
        product_shift[41]), .IN6(n67), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n53), .IN3(N106), .IN4(n68), .IN5(
        product_shift[40]), .IN6(n67), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n53), .IN3(N69), .IN4(n68), .IN5(
        product_shift[3]), .IN6(n67), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n53), .IN3(N105), .IN4(n68), .IN5(
        product_shift[39]), .IN6(n67), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n53), .IN3(N104), .IN4(n49), .IN5(
        product_shift[38]), .IN6(n46), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n53), .IN3(N103), .IN4(n48), .IN5(
        product_shift[37]), .IN6(n47), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n53), .IN3(N102), .IN4(n49), .IN5(
        product_shift[36]), .IN6(n46), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n53), .IN3(N101), .IN4(n48), .IN5(n3), .IN6(
        n47), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n53), .IN3(N100), .IN4(n49), .IN5(
        product_shift[34]), .IN6(n47), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n51), .IN3(N99), .IN4(n68), .IN5(n12), .IN6(
        n67), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n51), .IN3(N98), .IN4(n49), .IN5(n18), .IN6(
        n67), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n51), .IN3(N97), .IN4(n48), .IN5(n24), .IN6(
        n67), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n51), .IN3(N96), .IN4(n49), .IN5(n30), .IN6(
        n67), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n51), .IN3(N68), .IN4(n49), .IN5(
        product_shift[2]), .IN6(n67), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n51), .IN3(N95), .IN4(n49), .IN5(n36), .IN6(
        n67), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n51), .IN3(N94), .IN4(n49), .IN5(n42), .IN6(
        n67), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n51), .IN3(N93), .IN4(n49), .IN5(n44), .IN6(
        n67), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n51), .IN3(N92), .IN4(n49), .IN5(
        product_shift[26]), .IN6(n67), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n51), .IN3(N91), .IN4(n49), .IN5(
        product_shift[25]), .IN6(n67), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n51), .IN3(N90), .IN4(n49), .IN5(
        product_shift[24]), .IN6(n67), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n51), .IN3(N89), .IN4(n49), .IN5(
        product_shift[23]), .IN6(n67), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n52), .IN3(N88), .IN4(n48), .IN5(
        product_shift[22]), .IN6(n67), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n52), .IN3(N87), .IN4(n48), .IN5(
        product_shift[21]), .IN6(n46), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n52), .IN3(N86), .IN4(n48), .IN5(
        product_shift[20]), .IN6(n46), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n52), .IN3(N67), .IN4(n48), .IN5(n46), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n52), .IN3(N85), .IN4(n48), .IN5(
        product_shift[19]), .IN6(n46), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n52), .IN3(N84), .IN4(n48), .IN5(
        product_shift[18]), .IN6(n46), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n52), .IN3(N83), .IN4(n48), .IN5(
        product_shift[17]), .IN6(n46), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n52), .IN3(N82), .IN4(n48), .IN5(
        product_shift[16]), .IN6(n46), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n52), .IN3(N81), .IN4(n48), .IN5(
        product_shift[15]), .IN6(n46), .Q(product2[15]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n52), .IN3(N79), .IN4(n48), .IN5(
        product_shift[13]), .IN6(n46), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n52), .IN3(N78), .IN4(n48), .IN5(
        product_shift[12]), .IN6(n46), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n53), .IN3(N77), .IN4(n49), .IN5(
        product_shift[11]), .IN6(n46), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n53), .IN3(N76), .IN4(n49), .IN5(
        product_shift[10]), .IN6(n47), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n67) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n66), .Q(n68) );
  booth6_14_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], 
        n3, product_shift[34], n12, n18, n24, n30, n36, n42, n44, 
        product_shift[26:0]}), .B({combined_negative_b[24:8], n5, n14, n20, 
        n26, n32, n38, combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM({N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, 
        SYNOPSYS_UNCONNECTED__0, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, SYNOPSYS_UNCONNECTED__1}) );
  booth6_14_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n12, n18, n24, n30, n36, n42, n44, product_shift[26:0]}), .B({
        combined_b[24:8], n10, n16, n22, n28, n34, n40, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        SYNOPSYS_UNCONNECTED__2, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  NBUFFX2 U3 ( .INP(product_shift[35]), .Z(n3) );
  INVX0 U4 ( .INP(combined_negative_b[7]), .ZN(n4) );
  INVX0 U52 ( .INP(n4), .ZN(n5) );
  INVX0 U57 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U60 ( .INP(n9), .ZN(n10) );
  INVX0 U61 ( .INP(product_shift[33]), .ZN(n11) );
  INVX0 U62 ( .INP(n11), .ZN(n12) );
  INVX0 U63 ( .INP(combined_negative_b[6]), .ZN(n13) );
  INVX0 U64 ( .INP(n13), .ZN(n14) );
  INVX0 U65 ( .INP(combined_b[6]), .ZN(n15) );
  INVX0 U66 ( .INP(n15), .ZN(n16) );
  INVX0 U67 ( .INP(product_shift[32]), .ZN(n17) );
  INVX0 U68 ( .INP(n17), .ZN(n18) );
  INVX0 U69 ( .INP(combined_negative_b[5]), .ZN(n19) );
  INVX0 U70 ( .INP(n19), .ZN(n20) );
  INVX0 U71 ( .INP(combined_b[5]), .ZN(n21) );
  INVX0 U72 ( .INP(n21), .ZN(n22) );
  INVX0 U73 ( .INP(product_shift[31]), .ZN(n23) );
  INVX0 U74 ( .INP(n23), .ZN(n24) );
  INVX0 U75 ( .INP(combined_negative_b[4]), .ZN(n25) );
  INVX0 U76 ( .INP(n25), .ZN(n26) );
  INVX0 U77 ( .INP(combined_b[4]), .ZN(n27) );
  INVX0 U78 ( .INP(n27), .ZN(n28) );
  INVX0 U79 ( .INP(product_shift[30]), .ZN(n29) );
  INVX0 U80 ( .INP(n29), .ZN(n30) );
  INVX0 U81 ( .INP(combined_negative_b[3]), .ZN(n31) );
  INVX0 U82 ( .INP(n31), .ZN(n32) );
  INVX0 U83 ( .INP(combined_b[3]), .ZN(n33) );
  INVX0 U84 ( .INP(n33), .ZN(n34) );
  INVX0 U85 ( .INP(product_shift[29]), .ZN(n35) );
  INVX0 U86 ( .INP(n35), .ZN(n36) );
  INVX0 U87 ( .INP(combined_negative_b[2]), .ZN(n37) );
  INVX0 U88 ( .INP(n37), .ZN(n38) );
  INVX0 U89 ( .INP(combined_b[2]), .ZN(n39) );
  INVX0 U90 ( .INP(n39), .ZN(n40) );
  INVX0 U91 ( .INP(product_shift[28]), .ZN(n41) );
  INVX0 U92 ( .INP(n41), .ZN(n42) );
  NBUFFX2 U93 ( .INP(n45), .Z(n54) );
  NBUFFX2 U94 ( .INP(n45), .Z(n55) );
  NBUFFX2 U95 ( .INP(n45), .Z(n56) );
  NBUFFX2 U96 ( .INP(n45), .Z(n57) );
  NBUFFX2 U97 ( .INP(n45), .Z(n58) );
  NBUFFX2 U98 ( .INP(n45), .Z(n59) );
  NBUFFX2 U99 ( .INP(n45), .Z(n60) );
  NBUFFX2 U100 ( .INP(n45), .Z(n61) );
  NBUFFX2 U101 ( .INP(n45), .Z(n63) );
  NBUFFX2 U102 ( .INP(n45), .Z(n64) );
  NBUFFX2 U103 ( .INP(n45), .Z(n65) );
  NBUFFX2 U104 ( .INP(n45), .Z(n62) );
  NBUFFX2 U105 ( .INP(n69), .Z(n51) );
  NBUFFX2 U106 ( .INP(n69), .Z(n50) );
  NBUFFX2 U107 ( .INP(n69), .Z(n52) );
  NBUFFX2 U108 ( .INP(n69), .Z(n53) );
  NBUFFX2 U109 ( .INP(n67), .Z(n46) );
  NBUFFX2 U110 ( .INP(n67), .Z(n47) );
  NBUFFX2 U111 ( .INP(n68), .Z(n48) );
  NBUFFX2 U112 ( .INP(n68), .Z(n49) );
  NBUFFX2 U113 ( .INP(reset), .Z(n45) );
  NOR2X0 U114 ( .IN1(n66), .IN2(product_shift[1]), .QN(n69) );
  INVX0 U115 ( .INP(product_shift[0]), .ZN(n66) );
  INVX0 U117 ( .INP(product_shift[27]), .ZN(n43) );
  INVX0 U118 ( .INP(n43), .ZN(n44) );
endmodule


module booth6_13_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  XOR2X1 U2 ( .IN1(n16), .IN2(carry[41]), .Q(SUM[41]) );
  NAND3X0 U3 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(n12) );
  NAND3X0 U4 ( .IN1(n29), .IN2(n28), .IN3(n27), .QN(n11) );
  NAND2X0 U5 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U6 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U7 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U8 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U9 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U10 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U11 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U12 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U13 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U14 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XOR3X1 U15 ( .IN1(A[34]), .IN2(carry[34]), .IN3(B[34]), .Q(SUM[34]) );
  NAND2X1 U16 ( .IN1(B[34]), .IN2(A[34]), .QN(n8) );
  NAND2X1 U17 ( .IN1(carry[34]), .IN2(A[34]), .QN(n9) );
  NAND2X1 U18 ( .IN1(carry[34]), .IN2(B[34]), .QN(n10) );
  NAND3X0 U19 ( .IN1(n8), .IN2(n10), .IN3(n9), .QN(carry[35]) );
  AND2X1 U20 ( .IN1(A[26]), .IN2(B[26]), .Q(n37) );
  XOR3X1 U21 ( .IN1(B[27]), .IN2(n37), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U22 ( .IN1(n37), .IN2(B[27]), .QN(n35) );
  XOR3X1 U23 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X1 U24 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  XOR3X1 U25 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U26 ( .IN1(A[40]), .IN2(B[40]), .QN(n13) );
  NAND2X0 U27 ( .IN1(A[40]), .IN2(carry[40]), .QN(n14) );
  NAND2X0 U28 ( .IN1(B[40]), .IN2(carry[40]), .QN(n15) );
  NAND3X0 U29 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[41]) );
  XOR2X1 U30 ( .IN1(A[41]), .IN2(B[41]), .Q(n16) );
  NAND2X0 U31 ( .IN1(A[41]), .IN2(B[41]), .QN(n17) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(carry[41]), .QN(n18) );
  NAND2X0 U33 ( .IN1(B[41]), .IN2(carry[41]), .QN(n19) );
  NAND3X0 U34 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[42]) );
  NAND2X0 U35 ( .IN1(A[43]), .IN2(B[43]), .QN(n20) );
  NAND2X0 U36 ( .IN1(A[43]), .IN2(carry[43]), .QN(n21) );
  NAND2X0 U37 ( .IN1(B[43]), .IN2(carry[43]), .QN(n22) );
  NAND3X0 U38 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(carry[44]) );
  XOR2X1 U39 ( .IN1(A[44]), .IN2(B[44]), .Q(n23) );
  XOR2X1 U40 ( .IN1(n23), .IN2(n12), .Q(SUM[44]) );
  NAND2X0 U41 ( .IN1(A[44]), .IN2(B[44]), .QN(n24) );
  NAND2X0 U42 ( .IN1(A[44]), .IN2(carry[44]), .QN(n25) );
  NAND2X0 U43 ( .IN1(B[44]), .IN2(carry[44]), .QN(n26) );
  NAND3X0 U44 ( .IN1(n25), .IN2(n26), .IN3(n24), .QN(carry[45]) );
  NAND2X0 U45 ( .IN1(A[46]), .IN2(B[46]), .QN(n27) );
  NAND2X0 U46 ( .IN1(A[46]), .IN2(carry[46]), .QN(n28) );
  NAND2X0 U47 ( .IN1(B[46]), .IN2(carry[46]), .QN(n29) );
  NAND3X0 U48 ( .IN1(n29), .IN2(n28), .IN3(n27), .QN(carry[47]) );
  XOR2X1 U49 ( .IN1(A[47]), .IN2(B[47]), .Q(n30) );
  XOR2X1 U50 ( .IN1(n30), .IN2(n11), .Q(SUM[47]) );
  NAND2X0 U51 ( .IN1(A[47]), .IN2(B[47]), .QN(n31) );
  NAND2X0 U52 ( .IN1(A[47]), .IN2(carry[47]), .QN(n32) );
  NAND2X0 U53 ( .IN1(B[47]), .IN2(carry[47]), .QN(n33) );
  NAND3X0 U54 ( .IN1(n32), .IN2(n33), .IN3(n31), .QN(carry[48]) );
  NAND2X0 U55 ( .IN1(A[27]), .IN2(B[27]), .QN(n34) );
  NAND2X0 U56 ( .IN1(n37), .IN2(A[27]), .QN(n36) );
  NAND3X0 U57 ( .IN1(n34), .IN2(n36), .IN3(n35), .QN(carry[28]) );
  XOR2X1 U58 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_13_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n8), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR2X1 U6 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  XOR3X1 U7 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U8 ( .IN1(A[46]), .IN2(carry[46]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[46]), .IN2(carry[46]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[46]), .IN2(A[46]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[47]) );
  XOR3X1 U12 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  INVX0 U13 ( .INP(A[34]), .ZN(n7) );
  INVX0 U14 ( .INP(n7), .ZN(n8) );
  DELLN2X2 U15 ( .INP(carry[45]), .Z(n9) );
  XOR3X2 U16 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  AND2X1 U17 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  NAND2X0 U18 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  XOR3X2 U19 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U22 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U23 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U24 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U25 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U27 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U28 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U29 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[46]) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U32 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U33 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U34 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U40 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U41 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_13 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[13] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n73), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n73), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n16), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n22), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n28), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n34), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n40), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n5), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n14), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n20), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n26), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n32), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n38), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n65), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n65), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n64), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n62), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n62), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n62), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n62), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n62), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n62), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n62), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n62), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n62), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n62), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n57), .IN3(N75), .IN4(n52), .IN5(
        product_shift[9]), .IN6(n48), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n57), .IN3(N74), .IN4(n52), .IN5(
        product_shift[8]), .IN6(n51), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n57), .IN3(N73), .IN4(n52), .IN5(
        product_shift[7]), .IN6(n51), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n57), .IN3(N72), .IN4(n52), .IN5(
        product_shift[6]), .IN6(n51), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n57), .IN3(N71), .IN4(n52), .IN5(
        product_shift[5]), .IN6(n51), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n57), .IN3(N116), .IN4(n52), .IN5(
        product_shift[49]), .IN6(n51), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n57), .IN3(N70), .IN4(n52), .IN5(
        product_shift[4]), .IN6(n51), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n57), .IN3(N115), .IN4(n52), .IN5(
        product_shift[49]), .IN6(n51), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n57), .IN3(N114), .IN4(n52), .IN5(
        product_shift[48]), .IN6(n51), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n57), .IN3(N113), .IN4(n52), .IN5(
        product_shift[47]), .IN6(n51), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n57), .IN3(N112), .IN4(n52), .IN5(
        product_shift[46]), .IN6(n51), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n57), .IN3(N111), .IN4(n52), .IN5(
        product_shift[45]), .IN6(n51), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n58), .IN3(N110), .IN4(n53), .IN5(
        product_shift[44]), .IN6(n50), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n58), .IN3(N109), .IN4(n53), .IN5(
        product_shift[43]), .IN6(n50), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n58), .IN3(N108), .IN4(n53), .IN5(
        product_shift[42]), .IN6(n50), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n58), .IN3(N107), .IN4(n53), .IN5(
        product_shift[41]), .IN6(n50), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n58), .IN3(N106), .IN4(n53), .IN5(
        product_shift[40]), .IN6(n50), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n58), .IN3(N69), .IN4(n53), .IN5(
        product_shift[3]), .IN6(n50), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n58), .IN3(N105), .IN4(n53), .IN5(
        product_shift[39]), .IN6(n50), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n58), .IN3(N104), .IN4(n53), .IN5(
        product_shift[38]), .IN6(n50), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n58), .IN3(N103), .IN4(n53), .IN5(
        product_shift[37]), .IN6(n50), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n58), .IN3(N102), .IN4(n53), .IN5(
        product_shift[36]), .IN6(n50), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n58), .IN3(N101), .IN4(n53), .IN5(n3), .IN6(
        n50), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n58), .IN3(N100), .IN4(n53), .IN5(
        product_shift[34]), .IN6(n50), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n59), .IN3(N99), .IN4(n54), .IN5(n12), .IN6(
        n50), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n59), .IN3(N98), .IN4(n54), .IN5(n18), .IN6(
        n49), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n59), .IN3(N97), .IN4(n54), .IN5(n24), .IN6(
        n49), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n59), .IN3(N96), .IN4(n54), .IN5(n30), .IN6(
        n49), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n59), .IN3(N68), .IN4(n54), .IN5(
        product_shift[2]), .IN6(n49), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n59), .IN3(N95), .IN4(n54), .IN5(n36), .IN6(
        n49), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n59), .IN3(N94), .IN4(n54), .IN5(n42), .IN6(
        n49), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n59), .IN3(N93), .IN4(n54), .IN5(n44), .IN6(
        n49), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n59), .IN3(N92), .IN4(n54), .IN5(n46), .IN6(
        n49), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n59), .IN3(N91), .IN4(n54), .IN5(
        product_shift[25]), .IN6(n49), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n59), .IN3(N90), .IN4(n54), .IN5(
        product_shift[24]), .IN6(n49), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n59), .IN3(N89), .IN4(n54), .IN5(
        product_shift[23]), .IN6(n49), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n60), .IN3(N88), .IN4(n55), .IN5(
        product_shift[22]), .IN6(n49), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n60), .IN3(N87), .IN4(n55), .IN5(
        product_shift[21]), .IN6(n48), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n60), .IN3(N86), .IN4(n55), .IN5(
        product_shift[20]), .IN6(n48), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n60), .IN3(N67), .IN4(n55), .IN5(n48), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n60), .IN3(N85), .IN4(n55), .IN5(
        product_shift[19]), .IN6(n48), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n60), .IN3(N84), .IN4(n55), .IN5(
        product_shift[18]), .IN6(n48), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n60), .IN3(N83), .IN4(n55), .IN5(
        product_shift[17]), .IN6(n48), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n60), .IN3(N82), .IN4(n55), .IN5(
        product_shift[16]), .IN6(n48), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n60), .IN3(N81), .IN4(n55), .IN5(
        product_shift[15]), .IN6(n48), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n60), .IN3(N80), .IN4(n55), .IN5(
        product_shift[14]), .IN6(n48), .Q(product2[14]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n60), .IN3(N78), .IN4(n55), .IN5(
        product_shift[12]), .IN6(n48), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n61), .IN3(N77), .IN4(n56), .IN5(
        product_shift[11]), .IN6(n48), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n61), .IN3(N76), .IN4(n56), .IN5(
        product_shift[10]), .IN6(n49), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n75) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n74), .Q(n76) );
  booth6_13_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], 
        n3, product_shift[34], n12, n18, n24, n30, n36, n42, n44, n46, 
        product_shift[25:0]}), .B({combined_negative_b[24:8], n5, n14, n20, 
        n26, n32, n38, combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM({N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        SYNOPSYS_UNCONNECTED__0, N78, N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, SYNOPSYS_UNCONNECTED__1}) );
  booth6_13_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n12, n18, n24, n30, n36, n42, n44, n46, product_shift[25:0]}), .B({
        combined_b[24:8], n10, n16, n22, n28, n34, n40, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        SYNOPSYS_UNCONNECTED__2, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  NBUFFX2 U3 ( .INP(product_shift[35]), .Z(n3) );
  INVX0 U4 ( .INP(combined_negative_b[7]), .ZN(n4) );
  INVX0 U53 ( .INP(n4), .ZN(n5) );
  INVX0 U57 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U60 ( .INP(n9), .ZN(n10) );
  INVX0 U61 ( .INP(product_shift[33]), .ZN(n11) );
  INVX0 U62 ( .INP(n11), .ZN(n12) );
  INVX0 U63 ( .INP(combined_negative_b[6]), .ZN(n13) );
  INVX0 U64 ( .INP(n13), .ZN(n14) );
  INVX0 U65 ( .INP(combined_b[6]), .ZN(n15) );
  INVX0 U66 ( .INP(n15), .ZN(n16) );
  INVX0 U67 ( .INP(product_shift[32]), .ZN(n17) );
  INVX0 U68 ( .INP(n17), .ZN(n18) );
  INVX0 U69 ( .INP(combined_negative_b[5]), .ZN(n19) );
  INVX0 U70 ( .INP(n19), .ZN(n20) );
  INVX0 U71 ( .INP(combined_b[5]), .ZN(n21) );
  INVX0 U72 ( .INP(n21), .ZN(n22) );
  INVX0 U73 ( .INP(product_shift[31]), .ZN(n23) );
  INVX0 U74 ( .INP(n23), .ZN(n24) );
  INVX0 U75 ( .INP(combined_negative_b[4]), .ZN(n25) );
  INVX0 U76 ( .INP(n25), .ZN(n26) );
  INVX0 U77 ( .INP(combined_b[4]), .ZN(n27) );
  INVX0 U78 ( .INP(n27), .ZN(n28) );
  INVX0 U79 ( .INP(product_shift[30]), .ZN(n29) );
  INVX0 U80 ( .INP(n29), .ZN(n30) );
  INVX0 U81 ( .INP(combined_negative_b[3]), .ZN(n31) );
  INVX0 U82 ( .INP(n31), .ZN(n32) );
  INVX0 U83 ( .INP(combined_b[3]), .ZN(n33) );
  INVX0 U84 ( .INP(n33), .ZN(n34) );
  INVX0 U85 ( .INP(product_shift[29]), .ZN(n35) );
  INVX0 U86 ( .INP(n35), .ZN(n36) );
  INVX0 U87 ( .INP(combined_negative_b[2]), .ZN(n37) );
  INVX0 U88 ( .INP(n37), .ZN(n38) );
  INVX0 U89 ( .INP(combined_b[2]), .ZN(n39) );
  INVX0 U90 ( .INP(n39), .ZN(n40) );
  INVX0 U91 ( .INP(product_shift[28]), .ZN(n41) );
  INVX0 U92 ( .INP(n41), .ZN(n42) );
  NBUFFX2 U93 ( .INP(n47), .Z(n62) );
  NBUFFX2 U94 ( .INP(n47), .Z(n63) );
  NBUFFX2 U95 ( .INP(n47), .Z(n64) );
  NBUFFX2 U96 ( .INP(n47), .Z(n65) );
  NBUFFX2 U97 ( .INP(n47), .Z(n66) );
  NBUFFX2 U98 ( .INP(n47), .Z(n67) );
  NBUFFX2 U99 ( .INP(n47), .Z(n68) );
  NBUFFX2 U100 ( .INP(n47), .Z(n69) );
  NBUFFX2 U101 ( .INP(n47), .Z(n71) );
  NBUFFX2 U102 ( .INP(n47), .Z(n72) );
  NBUFFX2 U103 ( .INP(n47), .Z(n73) );
  NBUFFX2 U104 ( .INP(n47), .Z(n70) );
  NBUFFX2 U105 ( .INP(n77), .Z(n59) );
  NBUFFX2 U106 ( .INP(n77), .Z(n58) );
  NBUFFX2 U107 ( .INP(n77), .Z(n57) );
  NBUFFX2 U108 ( .INP(n77), .Z(n60) );
  NBUFFX2 U109 ( .INP(n77), .Z(n61) );
  NBUFFX2 U110 ( .INP(n75), .Z(n49) );
  NBUFFX2 U111 ( .INP(n75), .Z(n50) );
  NBUFFX2 U112 ( .INP(n75), .Z(n48) );
  NBUFFX2 U113 ( .INP(n75), .Z(n51) );
  NBUFFX2 U114 ( .INP(n76), .Z(n54) );
  NBUFFX2 U115 ( .INP(n76), .Z(n53) );
  NBUFFX2 U116 ( .INP(n76), .Z(n52) );
  NBUFFX2 U117 ( .INP(n76), .Z(n55) );
  NBUFFX2 U118 ( .INP(n76), .Z(n56) );
  NBUFFX2 U119 ( .INP(reset), .Z(n47) );
  NOR2X0 U120 ( .IN1(n74), .IN2(product_shift[1]), .QN(n77) );
  INVX0 U121 ( .INP(product_shift[0]), .ZN(n74) );
  INVX0 U123 ( .INP(product_shift[27]), .ZN(n43) );
  INVX0 U124 ( .INP(n43), .ZN(n44) );
  INVX0 U125 ( .INP(product_shift[26]), .ZN(n45) );
  INVX0 U126 ( .INP(n45), .ZN(n46) );
endmodule


module booth6_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X1 U1 ( .IN1(carry[45]), .IN2(B[45]), .IN3(A[45]), .Q(SUM[45]) );
  NAND2X0 U2 ( .IN1(A[45]), .IN2(carry[45]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[45]), .IN2(carry[45]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[45]), .IN2(A[45]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[46]) );
  XOR3X2 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U7 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U11 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U13 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  XOR3X2 U17 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  DELLN2X2 U18 ( .INP(carry[47]), .Z(n11) );
  DELLN2X2 U19 ( .INP(carry[41]), .Z(n12) );
  DELLN2X2 U20 ( .INP(carry[44]), .Z(n13) );
  AND2X1 U21 ( .IN1(A[26]), .IN2(B[26]), .Q(n38) );
  XOR3X1 U22 ( .IN1(B[27]), .IN2(n38), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U23 ( .IN1(n38), .IN2(B[27]), .QN(n36) );
  XOR3X1 U24 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X1 U25 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U26 ( .IN1(A[40]), .IN2(B[40]), .QN(n14) );
  NAND2X0 U27 ( .IN1(A[40]), .IN2(carry[40]), .QN(n15) );
  NAND2X0 U28 ( .IN1(B[40]), .IN2(carry[40]), .QN(n16) );
  NAND3X0 U29 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(carry[41]) );
  XOR2X1 U30 ( .IN1(A[41]), .IN2(B[41]), .Q(n17) );
  XOR2X1 U31 ( .IN1(n17), .IN2(n12), .Q(SUM[41]) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(B[41]), .QN(n18) );
  NAND2X0 U33 ( .IN1(A[41]), .IN2(carry[41]), .QN(n19) );
  NAND2X0 U34 ( .IN1(B[41]), .IN2(carry[41]), .QN(n20) );
  NAND3X0 U35 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[42]) );
  NAND2X0 U36 ( .IN1(A[43]), .IN2(B[43]), .QN(n21) );
  NAND2X0 U37 ( .IN1(A[43]), .IN2(carry[43]), .QN(n22) );
  NAND2X0 U38 ( .IN1(B[43]), .IN2(carry[43]), .QN(n23) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n23), .IN3(n21), .QN(carry[44]) );
  XOR2X1 U40 ( .IN1(A[44]), .IN2(B[44]), .Q(n24) );
  XOR2X1 U41 ( .IN1(n24), .IN2(n13), .Q(SUM[44]) );
  NAND2X0 U42 ( .IN1(A[44]), .IN2(B[44]), .QN(n25) );
  NAND2X0 U43 ( .IN1(A[44]), .IN2(carry[44]), .QN(n26) );
  NAND2X0 U44 ( .IN1(B[44]), .IN2(carry[44]), .QN(n27) );
  NAND3X0 U45 ( .IN1(n26), .IN2(n27), .IN3(n25), .QN(carry[45]) );
  NAND2X0 U46 ( .IN1(A[46]), .IN2(B[46]), .QN(n28) );
  NAND2X0 U47 ( .IN1(A[46]), .IN2(carry[46]), .QN(n29) );
  NAND2X0 U48 ( .IN1(B[46]), .IN2(carry[46]), .QN(n30) );
  NAND3X0 U49 ( .IN1(n29), .IN2(n30), .IN3(n28), .QN(carry[47]) );
  XOR2X1 U50 ( .IN1(A[47]), .IN2(B[47]), .Q(n31) );
  XOR2X1 U51 ( .IN1(n31), .IN2(n11), .Q(SUM[47]) );
  NAND2X0 U52 ( .IN1(A[47]), .IN2(B[47]), .QN(n32) );
  NAND2X0 U53 ( .IN1(A[47]), .IN2(carry[47]), .QN(n33) );
  NAND2X0 U54 ( .IN1(B[47]), .IN2(carry[47]), .QN(n34) );
  NAND3X0 U55 ( .IN1(n33), .IN2(n34), .IN3(n32), .QN(carry[48]) );
  NAND2X0 U56 ( .IN1(A[27]), .IN2(B[27]), .QN(n35) );
  NAND2X0 U57 ( .IN1(n38), .IN2(A[27]), .QN(n37) );
  NAND3X0 U58 ( .IN1(n35), .IN2(n37), .IN3(n36), .QN(carry[28]) );
  XOR2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_12_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX2 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX2 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX2 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX2 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  XOR3X1 U1 ( .IN1(A[37]), .IN2(B[37]), .IN3(carry[37]), .Q(SUM[37]) );
  NAND2X0 U2 ( .IN1(A[37]), .IN2(B[37]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[37]), .IN2(carry[37]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[37]), .IN2(carry[37]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[38]) );
  XOR2X1 U6 ( .IN1(A[38]), .IN2(B[38]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[38]), .Q(SUM[38]) );
  NAND2X0 U8 ( .IN1(A[38]), .IN2(B[38]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[38]), .IN2(carry[38]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[38]), .IN2(carry[38]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[39]) );
  XOR2X1 U12 ( .IN1(n21), .IN2(carry[48]), .Q(SUM[48]) );
  XOR3X1 U13 ( .IN1(B[27]), .IN2(n28), .IN3(A[27]), .Q(SUM[27]) );
  INVX0 U14 ( .INP(A[34]), .ZN(n8) );
  INVX0 U15 ( .INP(n8), .ZN(n9) );
  DELLN2X2 U16 ( .INP(carry[45]), .Z(n10) );
  XOR3X2 U17 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  AND2X1 U18 ( .IN1(A[26]), .IN2(B[26]), .Q(n28) );
  NAND2X0 U19 ( .IN1(n28), .IN2(B[27]), .QN(n26) );
  XOR3X2 U20 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(B[44]), .QN(n11) );
  NAND2X0 U22 ( .IN1(A[44]), .IN2(carry[44]), .QN(n12) );
  NAND2X0 U23 ( .IN1(B[44]), .IN2(carry[44]), .QN(n13) );
  NAND3X0 U24 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[45]) );
  XOR2X1 U25 ( .IN1(A[45]), .IN2(B[45]), .Q(n14) );
  XOR2X1 U26 ( .IN1(n14), .IN2(n10), .Q(SUM[45]) );
  NAND2X0 U27 ( .IN1(A[45]), .IN2(B[45]), .QN(n15) );
  NAND2X0 U28 ( .IN1(A[45]), .IN2(carry[45]), .QN(n16) );
  NAND2X0 U29 ( .IN1(B[45]), .IN2(carry[45]), .QN(n17) );
  NAND3X0 U30 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[46]) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(B[47]), .QN(n18) );
  NAND2X0 U32 ( .IN1(A[47]), .IN2(carry[47]), .QN(n19) );
  NAND2X0 U33 ( .IN1(B[47]), .IN2(carry[47]), .QN(n20) );
  NAND3X0 U34 ( .IN1(n20), .IN2(n19), .IN3(n18), .QN(carry[48]) );
  XOR2X1 U35 ( .IN1(A[48]), .IN2(B[48]), .Q(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(B[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(A[48]), .IN2(carry[48]), .QN(n23) );
  NAND2X0 U38 ( .IN1(B[48]), .IN2(carry[48]), .QN(n24) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[49]) );
  NAND2X0 U40 ( .IN1(A[27]), .IN2(B[27]), .QN(n25) );
  NAND2X0 U41 ( .IN1(n28), .IN2(A[27]), .QN(n27) );
  NAND3X0 U42 ( .IN1(n25), .IN2(n27), .IN3(n26), .QN(carry[28]) );
  XOR2X1 U43 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_12 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[12] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n73), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n73), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n68), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n16), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n22), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n28), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n34), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n40), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n67), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n66), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n5), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n14), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n20), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n26), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n32), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n38), .CLK(clk), .RSTB(n65), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n65), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n65), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n64), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n64), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n62), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n62), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n62), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n62), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n62), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n62), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n62), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n62), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n62), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n62), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n62), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n57), .IN3(N75), .IN4(n52), .IN5(
        product_shift[9]), .IN6(n48), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n57), .IN3(N74), .IN4(n52), .IN5(
        product_shift[8]), .IN6(n51), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n57), .IN3(N73), .IN4(n52), .IN5(
        product_shift[7]), .IN6(n51), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n57), .IN3(N72), .IN4(n52), .IN5(
        product_shift[6]), .IN6(n51), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n57), .IN3(N71), .IN4(n52), .IN5(
        product_shift[5]), .IN6(n51), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n57), .IN3(N116), .IN4(n52), .IN5(
        product_shift[49]), .IN6(n51), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n57), .IN3(N70), .IN4(n52), .IN5(
        product_shift[4]), .IN6(n51), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n57), .IN3(N115), .IN4(n52), .IN5(
        product_shift[49]), .IN6(n51), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n57), .IN3(N114), .IN4(n52), .IN5(
        product_shift[48]), .IN6(n51), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n57), .IN3(N113), .IN4(n52), .IN5(
        product_shift[47]), .IN6(n51), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n57), .IN3(N112), .IN4(n52), .IN5(
        product_shift[46]), .IN6(n51), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n57), .IN3(N111), .IN4(n52), .IN5(
        product_shift[45]), .IN6(n51), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n58), .IN3(N110), .IN4(n53), .IN5(
        product_shift[44]), .IN6(n50), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n58), .IN3(N109), .IN4(n53), .IN5(
        product_shift[43]), .IN6(n50), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n58), .IN3(N108), .IN4(n53), .IN5(
        product_shift[42]), .IN6(n50), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n58), .IN3(N107), .IN4(n53), .IN5(
        product_shift[41]), .IN6(n50), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n58), .IN3(N106), .IN4(n53), .IN5(
        product_shift[40]), .IN6(n50), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n58), .IN3(N69), .IN4(n53), .IN5(
        product_shift[3]), .IN6(n50), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n58), .IN3(N105), .IN4(n53), .IN5(
        product_shift[39]), .IN6(n50), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n58), .IN3(N104), .IN4(n53), .IN5(
        product_shift[38]), .IN6(n50), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n58), .IN3(N103), .IN4(n53), .IN5(
        product_shift[37]), .IN6(n50), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n58), .IN3(N102), .IN4(n53), .IN5(
        product_shift[36]), .IN6(n50), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n58), .IN3(N101), .IN4(n53), .IN5(n3), .IN6(
        n50), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n58), .IN3(N100), .IN4(n53), .IN5(
        product_shift[34]), .IN6(n50), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n59), .IN3(N99), .IN4(n54), .IN5(n12), .IN6(
        n50), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n59), .IN3(N98), .IN4(n54), .IN5(n18), .IN6(
        n49), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n59), .IN3(N97), .IN4(n54), .IN5(n24), .IN6(
        n49), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n59), .IN3(N96), .IN4(n54), .IN5(n30), .IN6(
        n49), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n59), .IN3(N68), .IN4(n54), .IN5(
        product_shift[2]), .IN6(n49), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n59), .IN3(N95), .IN4(n54), .IN5(n36), .IN6(
        n49), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n59), .IN3(N94), .IN4(n54), .IN5(n42), .IN6(
        n49), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n59), .IN3(N93), .IN4(n54), .IN5(n44), .IN6(
        n49), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n59), .IN3(N92), .IN4(n54), .IN5(n46), .IN6(
        n49), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n59), .IN3(N91), .IN4(n54), .IN5(
        product_shift[25]), .IN6(n49), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n59), .IN3(N90), .IN4(n54), .IN5(
        product_shift[24]), .IN6(n49), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n59), .IN3(N89), .IN4(n54), .IN5(
        product_shift[23]), .IN6(n49), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n60), .IN3(N88), .IN4(n55), .IN5(
        product_shift[22]), .IN6(n49), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n60), .IN3(N87), .IN4(n55), .IN5(
        product_shift[21]), .IN6(n48), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n60), .IN3(N86), .IN4(n55), .IN5(
        product_shift[20]), .IN6(n48), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n60), .IN3(N67), .IN4(n55), .IN5(n48), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n60), .IN3(N85), .IN4(n55), .IN5(
        product_shift[19]), .IN6(n48), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n60), .IN3(N84), .IN4(n55), .IN5(
        product_shift[18]), .IN6(n48), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n60), .IN3(N83), .IN4(n55), .IN5(
        product_shift[17]), .IN6(n48), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n60), .IN3(N82), .IN4(n55), .IN5(
        product_shift[16]), .IN6(n48), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n60), .IN3(N81), .IN4(n55), .IN5(
        product_shift[15]), .IN6(n48), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n60), .IN3(N80), .IN4(n55), .IN5(
        product_shift[14]), .IN6(n48), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n60), .IN3(N79), .IN4(n55), .IN5(
        product_shift[13]), .IN6(n48), .Q(product2[13]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n61), .IN3(N77), .IN4(n56), .IN5(
        product_shift[11]), .IN6(n48), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n61), .IN3(N76), .IN4(n56), .IN5(
        product_shift[10]), .IN6(n49), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n75) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n74), .Q(n76) );
  booth6_12_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], 
        n3, product_shift[34], n12, n18, n24, n30, n36, n42, n44, n46, 
        product_shift[25:0]}), .B({combined_negative_b[24:8], n5, n14, n20, 
        n26, n32, n38, combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM({N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        SYNOPSYS_UNCONNECTED__0, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, SYNOPSYS_UNCONNECTED__1}) );
  booth6_12_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n12, n18, n24, n30, n36, n42, n44, n46, product_shift[25:0]}), .B({
        combined_b[24:8], n10, n16, n22, n28, n34, n40, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, SYNOPSYS_UNCONNECTED__2, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n47), .Q(
        product2_o[36]) );
  NBUFFX2 U3 ( .INP(product_shift[35]), .Z(n3) );
  INVX0 U4 ( .INP(combined_negative_b[7]), .ZN(n4) );
  INVX0 U54 ( .INP(n4), .ZN(n5) );
  INVX0 U57 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U60 ( .INP(n9), .ZN(n10) );
  INVX0 U61 ( .INP(product_shift[33]), .ZN(n11) );
  INVX0 U62 ( .INP(n11), .ZN(n12) );
  INVX0 U63 ( .INP(combined_negative_b[6]), .ZN(n13) );
  INVX0 U64 ( .INP(n13), .ZN(n14) );
  INVX0 U65 ( .INP(combined_b[6]), .ZN(n15) );
  INVX0 U66 ( .INP(n15), .ZN(n16) );
  INVX0 U67 ( .INP(product_shift[32]), .ZN(n17) );
  INVX0 U68 ( .INP(n17), .ZN(n18) );
  INVX0 U69 ( .INP(combined_negative_b[5]), .ZN(n19) );
  INVX0 U70 ( .INP(n19), .ZN(n20) );
  INVX0 U71 ( .INP(combined_b[5]), .ZN(n21) );
  INVX0 U72 ( .INP(n21), .ZN(n22) );
  INVX0 U73 ( .INP(product_shift[31]), .ZN(n23) );
  INVX0 U74 ( .INP(n23), .ZN(n24) );
  INVX0 U75 ( .INP(combined_negative_b[4]), .ZN(n25) );
  INVX0 U76 ( .INP(n25), .ZN(n26) );
  INVX0 U77 ( .INP(combined_b[4]), .ZN(n27) );
  INVX0 U78 ( .INP(n27), .ZN(n28) );
  INVX0 U79 ( .INP(product_shift[30]), .ZN(n29) );
  INVX0 U80 ( .INP(n29), .ZN(n30) );
  INVX0 U81 ( .INP(combined_negative_b[3]), .ZN(n31) );
  INVX0 U82 ( .INP(n31), .ZN(n32) );
  INVX0 U83 ( .INP(combined_b[3]), .ZN(n33) );
  INVX0 U84 ( .INP(n33), .ZN(n34) );
  INVX0 U85 ( .INP(product_shift[29]), .ZN(n35) );
  INVX0 U86 ( .INP(n35), .ZN(n36) );
  INVX0 U87 ( .INP(combined_negative_b[2]), .ZN(n37) );
  INVX0 U88 ( .INP(n37), .ZN(n38) );
  INVX0 U89 ( .INP(combined_b[2]), .ZN(n39) );
  INVX0 U90 ( .INP(n39), .ZN(n40) );
  INVX0 U91 ( .INP(product_shift[28]), .ZN(n41) );
  INVX0 U92 ( .INP(n41), .ZN(n42) );
  NBUFFX2 U93 ( .INP(n47), .Z(n62) );
  NBUFFX2 U94 ( .INP(n72), .Z(n63) );
  NBUFFX2 U95 ( .INP(n47), .Z(n64) );
  NBUFFX2 U96 ( .INP(n70), .Z(n65) );
  NBUFFX2 U97 ( .INP(n47), .Z(n66) );
  NBUFFX2 U98 ( .INP(n47), .Z(n67) );
  NBUFFX2 U99 ( .INP(n47), .Z(n68) );
  NBUFFX2 U100 ( .INP(n47), .Z(n69) );
  NBUFFX2 U101 ( .INP(n47), .Z(n71) );
  NBUFFX2 U102 ( .INP(n47), .Z(n72) );
  NBUFFX2 U103 ( .INP(n47), .Z(n73) );
  NBUFFX2 U104 ( .INP(n47), .Z(n70) );
  NBUFFX2 U105 ( .INP(n77), .Z(n59) );
  NBUFFX2 U106 ( .INP(n77), .Z(n58) );
  NBUFFX2 U107 ( .INP(n77), .Z(n57) );
  NBUFFX2 U108 ( .INP(n77), .Z(n60) );
  NBUFFX2 U109 ( .INP(n77), .Z(n61) );
  NBUFFX2 U110 ( .INP(n75), .Z(n49) );
  NBUFFX2 U111 ( .INP(n75), .Z(n50) );
  NBUFFX2 U112 ( .INP(n75), .Z(n48) );
  NBUFFX2 U113 ( .INP(n75), .Z(n51) );
  NBUFFX2 U114 ( .INP(n76), .Z(n54) );
  NBUFFX2 U115 ( .INP(n76), .Z(n53) );
  NBUFFX2 U116 ( .INP(n76), .Z(n52) );
  NBUFFX2 U117 ( .INP(n76), .Z(n55) );
  NBUFFX2 U118 ( .INP(n76), .Z(n56) );
  NBUFFX2 U119 ( .INP(reset), .Z(n47) );
  NOR2X0 U120 ( .IN1(n74), .IN2(product_shift[1]), .QN(n77) );
  INVX0 U121 ( .INP(product_shift[0]), .ZN(n74) );
  INVX0 U123 ( .INP(product_shift[27]), .ZN(n43) );
  INVX0 U124 ( .INP(n43), .ZN(n44) );
  INVX0 U125 ( .INP(product_shift[26]), .ZN(n45) );
  INVX0 U126 ( .INP(n45), .ZN(n46) );
endmodule


module booth6_11_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   \carry[50] , \carry[49] , \carry[48] , \carry[47] , \carry[46] ,
         \carry[45] , \carry[44] , \carry[43] , \carry[42] , \carry[41] ,
         \carry[40] , \carry[39] , \carry[38] , \carry[37] , \carry[36] ,
         \carry[35] , \carry[34] , \carry[33] , \carry[32] , \carry[31] ,
         \carry[30] , \carry[29] , \carry[28] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n32), .CO(\carry[28] ), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(\carry[50] ), .Q(SUM[50]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(\carry[36] ), .CO(\carry[37] ), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(\carry[34] ), .CO(\carry[35] ), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(\carry[33] ), .CO(\carry[34] ), .S(
        SUM[33]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(\carry[45] ), .CO(\carry[46] ), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(\carry[44] ), .CO(\carry[45] ), .S(
        SUM[44]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(\carry[39] ), .CO(\carry[40] ), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(\carry[38] ), .CO(\carry[39] ), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(\carry[37] ), .CO(\carry[38] ), .S(
        SUM[37]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(\carry[47] ), .CO(\carry[48] ), .S(
        SUM[47]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(\carry[46] ), .CO(\carry[47] ), .S(
        SUM[46]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(\carry[41] ), .CO(\carry[42] ), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(\carry[40] ), .CO(\carry[41] ), .S(
        SUM[40]) );
  XOR3X1 U1 ( .IN1(A[29]), .IN2(B[29]), .IN3(\carry[29] ), .Q(SUM[29]) );
  XOR2X1 U2 ( .IN1(A[30]), .IN2(B[30]), .Q(n25) );
  XOR3X1 U3 ( .IN1(A[31]), .IN2(B[31]), .IN3(\carry[31] ), .Q(SUM[31]) );
  XOR2X1 U4 ( .IN1(A[32]), .IN2(B[32]), .Q(n18) );
  XOR3X1 U5 ( .IN1(A[42]), .IN2(B[42]), .IN3(\carry[42] ), .Q(SUM[42]) );
  XOR3X1 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(\carry[48] ), .Q(SUM[48]) );
  NAND2X0 U7 ( .IN1(A[48]), .IN2(B[48]), .QN(n1) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(\carry[48] ), .QN(n2) );
  NAND2X0 U9 ( .IN1(B[48]), .IN2(\carry[48] ), .QN(n3) );
  NAND3X0 U10 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(\carry[49] ) );
  XOR2X1 U11 ( .IN1(A[49]), .IN2(B[49]), .Q(n4) );
  XOR2X1 U12 ( .IN1(n4), .IN2(\carry[49] ), .Q(SUM[49]) );
  NAND2X0 U13 ( .IN1(A[49]), .IN2(B[49]), .QN(n5) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(\carry[49] ), .QN(n6) );
  NAND2X0 U15 ( .IN1(B[49]), .IN2(\carry[49] ), .QN(n7) );
  NAND3X0 U16 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(\carry[50] ) );
  NAND2X0 U17 ( .IN1(A[42]), .IN2(B[42]), .QN(n8) );
  NAND2X0 U18 ( .IN1(A[42]), .IN2(\carry[42] ), .QN(n9) );
  NAND2X0 U19 ( .IN1(B[42]), .IN2(\carry[42] ), .QN(n10) );
  NAND3X0 U20 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(\carry[43] ) );
  XOR2X1 U21 ( .IN1(A[43]), .IN2(B[43]), .Q(n11) );
  XOR2X1 U22 ( .IN1(n11), .IN2(\carry[43] ), .Q(SUM[43]) );
  NAND2X0 U23 ( .IN1(A[43]), .IN2(B[43]), .QN(n12) );
  NAND2X0 U24 ( .IN1(A[43]), .IN2(\carry[43] ), .QN(n13) );
  NAND2X0 U25 ( .IN1(B[43]), .IN2(\carry[43] ), .QN(n14) );
  NAND3X0 U26 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(\carry[44] ) );
  NAND2X0 U27 ( .IN1(A[31]), .IN2(B[31]), .QN(n15) );
  NAND2X0 U28 ( .IN1(A[31]), .IN2(\carry[31] ), .QN(n16) );
  NAND2X0 U29 ( .IN1(B[31]), .IN2(\carry[31] ), .QN(n17) );
  NAND3X0 U30 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(\carry[32] ) );
  XOR2X1 U31 ( .IN1(n18), .IN2(\carry[32] ), .Q(SUM[32]) );
  NAND2X0 U32 ( .IN1(A[32]), .IN2(B[32]), .QN(n19) );
  NAND2X0 U33 ( .IN1(A[32]), .IN2(\carry[32] ), .QN(n20) );
  NAND2X0 U34 ( .IN1(B[32]), .IN2(\carry[32] ), .QN(n21) );
  NAND3X0 U35 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(\carry[33] ) );
  NAND2X0 U36 ( .IN1(A[29]), .IN2(B[29]), .QN(n22) );
  NAND2X0 U37 ( .IN1(A[29]), .IN2(\carry[29] ), .QN(n23) );
  NAND2X0 U38 ( .IN1(B[29]), .IN2(\carry[29] ), .QN(n24) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(\carry[30] ) );
  XOR2X1 U40 ( .IN1(n25), .IN2(\carry[30] ), .Q(SUM[30]) );
  NAND2X0 U41 ( .IN1(A[30]), .IN2(B[30]), .QN(n26) );
  NAND2X0 U42 ( .IN1(A[30]), .IN2(\carry[30] ), .QN(n27) );
  NAND2X0 U43 ( .IN1(B[30]), .IN2(\carry[30] ), .QN(n28) );
  NAND3X0 U44 ( .IN1(n26), .IN2(n27), .IN3(n28), .QN(\carry[31] ) );
  XOR3X1 U45 ( .IN1(\carry[35] ), .IN2(A[35]), .IN3(B[35]), .Q(SUM[35]) );
  NAND2X0 U46 ( .IN1(B[35]), .IN2(\carry[35] ), .QN(n29) );
  NAND2X0 U47 ( .IN1(A[35]), .IN2(\carry[35] ), .QN(n30) );
  NAND2X0 U48 ( .IN1(A[35]), .IN2(B[35]), .QN(n31) );
  NAND3X0 U49 ( .IN1(n29), .IN2(n31), .IN3(n30), .QN(\carry[36] ) );
  AND2X1 U50 ( .IN1(A[26]), .IN2(B[26]), .Q(n32) );
  XOR2X1 U51 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_11_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X1 U1 ( .IN1(carry[41]), .IN2(B[41]), .IN3(A[41]), .Q(SUM[41]) );
  NAND2X1 U2 ( .IN1(A[41]), .IN2(carry[41]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[41]), .IN2(carry[41]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[41]), .IN2(A[41]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[42]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n26), .IN3(A[27]), .Q(SUM[27]) );
  XNOR2X1 U7 ( .IN1(n19), .IN2(n7), .Q(SUM[48]) );
  XOR3X1 U8 ( .IN1(B[35]), .IN2(A[35]), .IN3(carry[35]), .Q(SUM[35]) );
  NAND2X1 U9 ( .IN1(carry[35]), .IN2(B[35]), .QN(n4) );
  NAND2X1 U10 ( .IN1(A[35]), .IN2(B[35]), .QN(n5) );
  NAND2X0 U11 ( .IN1(A[35]), .IN2(carry[35]), .QN(n6) );
  NAND3X0 U12 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[36]) );
  INVX0 U13 ( .INP(carry[48]), .ZN(n7) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n8) );
  XOR3X2 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  AND2X1 U16 ( .IN1(A[26]), .IN2(B[26]), .Q(n26) );
  NAND2X0 U17 ( .IN1(n26), .IN2(B[27]), .QN(n24) );
  XOR3X2 U18 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n9) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n10) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n11) );
  NAND3X0 U22 ( .IN1(n11), .IN2(n10), .IN3(n9), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n12) );
  XOR2X1 U24 ( .IN1(n12), .IN2(n8), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n13) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n14) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n15) );
  NAND3X0 U28 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[46]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n16) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n17) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n18) );
  NAND3X0 U32 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n19) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(B[48]), .QN(n20) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(carry[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(B[48]), .IN2(carry[48]), .QN(n22) );
  NAND3X0 U37 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(carry[49]) );
  NAND2X0 U38 ( .IN1(A[27]), .IN2(B[27]), .QN(n23) );
  NAND2X0 U39 ( .IN1(n26), .IN2(A[27]), .QN(n25) );
  NAND3X0 U40 ( .IN1(n23), .IN2(n25), .IN3(n24), .QN(carry[28]) );
  XOR2X1 U41 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_11 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n6, n7, net20870, net20868, net20866,
         net20864, net20876, net20874, net20888, net20886, n3, n4, n5, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[11] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n67), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n67), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n63), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n62), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n62), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n10), .CLK(clk), .RSTB(n62), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n16), .CLK(clk), .RSTB(n62), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n22), .CLK(clk), .RSTB(n62), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n28), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n34), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n40), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n61), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n60), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n12), .CLK(clk), .RSTB(n60), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n18), .CLK(clk), .RSTB(n60), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n24), .CLK(clk), .RSTB(n60), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n30), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n36), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n42), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n46), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n50), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n59), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n58), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n56), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n56), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n56), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n56), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n56), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n56), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n56), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n56), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n56), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n56), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(net20864), .IN3(N75), .IN4(net20874), .IN5(
        product_shift[9]), .IN6(n5), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(net20864), .IN3(N74), .IN4(net20874), .IN5(
        product_shift[8]), .IN6(net20886), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(net20864), .IN3(N73), .IN4(net20874), .IN5(
        product_shift[7]), .IN6(net20888), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(net20864), .IN3(N72), .IN4(net20874), .IN5(
        product_shift[6]), .IN6(n5), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(net20864), .IN3(N71), .IN4(net20874), .IN5(
        product_shift[5]), .IN6(n5), .Q(product2[5]) );
  AO222X1 U13 ( .IN1(N19), .IN2(net20864), .IN3(N70), .IN4(net20874), .IN5(
        product_shift[4]), .IN6(n5), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(net20864), .IN3(N115), .IN4(net20874), .IN5(
        product_shift[49]), .IN6(n5), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(net20864), .IN3(N114), .IN4(net20874), .IN5(
        product_shift[48]), .IN6(n5), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(net20864), .IN3(N113), .IN4(net20874), .IN5(
        product_shift[47]), .IN6(n5), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(net20864), .IN3(N112), .IN4(net20874), .IN5(
        product_shift[46]), .IN6(n5), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(net20864), .IN3(N111), .IN4(net20874), .IN5(
        product_shift[45]), .IN6(n5), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(net20866), .IN3(N110), .IN4(net20876), .IN5(
        product_shift[44]), .IN6(net20888), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(net20866), .IN3(N109), .IN4(net20876), .IN5(
        product_shift[43]), .IN6(net20888), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(net20866), .IN3(N108), .IN4(net20876), .IN5(
        product_shift[42]), .IN6(net20888), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(net20866), .IN3(N107), .IN4(net20876), .IN5(
        product_shift[41]), .IN6(net20888), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(net20866), .IN3(N106), .IN4(net20876), .IN5(
        product_shift[40]), .IN6(net20888), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(net20866), .IN3(N69), .IN4(net20876), .IN5(
        product_shift[3]), .IN6(net20888), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(net20866), .IN3(N105), .IN4(net20876), .IN5(
        product_shift[39]), .IN6(net20888), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(net20866), .IN3(N104), .IN4(net20876), .IN5(
        product_shift[38]), .IN6(net20888), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(net20866), .IN3(N103), .IN4(net20876), .IN5(
        product_shift[37]), .IN6(net20888), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(net20866), .IN3(N102), .IN4(net20876), .IN5(
        product_shift[36]), .IN6(net20888), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(net20866), .IN3(N101), .IN4(net20876), .IN5(n4), .IN6(net20888), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(net20866), .IN3(N100), .IN4(net20876), .IN5(
        n14), .IN6(net20888), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(net20868), .IN3(N99), .IN4(n7), .IN5(n20), 
        .IN6(net20888), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(net20868), .IN3(N98), .IN4(net20876), .IN5(n26), .IN6(net20886), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(net20868), .IN3(N97), .IN4(net20874), .IN5(n32), .IN6(net20886), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(net20868), .IN3(N96), .IN4(net20876), .IN5(n38), .IN6(net20886), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(net20868), .IN3(N68), .IN4(n7), .IN5(
        product_shift[2]), .IN6(net20886), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(net20868), .IN3(N95), .IN4(n7), .IN5(n44), 
        .IN6(net20886), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(net20868), .IN3(N94), .IN4(n7), .IN5(n48), 
        .IN6(net20886), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(net20868), .IN3(N93), .IN4(n7), .IN5(n52), 
        .IN6(net20886), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(net20868), .IN3(N92), .IN4(n7), .IN5(n54), 
        .IN6(net20886), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(net20868), .IN3(N91), .IN4(n7), .IN5(
        product_shift[25]), .IN6(net20886), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(net20868), .IN3(N90), .IN4(n7), .IN5(
        product_shift[24]), .IN6(net20886), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(net20868), .IN3(N89), .IN4(n7), .IN5(
        product_shift[23]), .IN6(net20886), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(net20870), .IN3(N88), .IN4(n7), .IN5(
        product_shift[22]), .IN6(net20886), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(net20870), .IN3(N87), .IN4(n7), .IN5(
        product_shift[21]), .IN6(net20886), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(net20870), .IN3(N86), .IN4(n7), .IN5(
        product_shift[20]), .IN6(net20888), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(net20870), .IN3(N67), .IN4(net20874), .IN5(n5), 
        .IN6(product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(net20870), .IN3(N85), .IN4(n7), .IN5(
        product_shift[19]), .IN6(n5), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(net20870), .IN3(N84), .IN4(n7), .IN5(
        product_shift[18]), .IN6(n5), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(net20870), .IN3(N83), .IN4(n7), .IN5(
        product_shift[17]), .IN6(n5), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(net20870), .IN3(N82), .IN4(n7), .IN5(
        product_shift[16]), .IN6(n5), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(net20870), .IN3(N81), .IN4(n7), .IN5(
        product_shift[15]), .IN6(n5), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(net20870), .IN3(N80), .IN4(n7), .IN5(
        product_shift[14]), .IN6(n5), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(net20870), .IN3(N79), .IN4(n7), .IN5(
        product_shift[13]), .IN6(n5), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(net20870), .IN3(N78), .IN4(n7), .IN5(
        product_shift[12]), .IN6(n5), .Q(product2[12]) );
  AO222X1 U56 ( .IN1(N25), .IN2(net20870), .IN3(N76), .IN4(net20876), .IN5(
        product_shift[10]), .IN6(net20886), .Q(product2[10]) );
  booth6_11_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], 
        n4, n14, n20, n26, n32, n38, n44, n48, n52, n54, product_shift[25:0]}), 
        .B({combined_negative_b[24:9], n12, n18, n24, n30, n36, n42, n46, n50, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, 
        SYNOPSYS_UNCONNECTED__0, N76, N75, N74, N73, N72, N71, N70, N69, N68, 
        N67, SYNOPSYS_UNCONNECTED__1}) );
  booth6_11_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:36], 
        n4, n14, n20, n26, n32, n38, n44, n48, n52, n54, product_shift[25:0]}), 
        .B({combined_b[24:8], n10, n16, n22, n28, n34, n40, combined_b[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, SYNOPSYS_UNCONNECTED__2, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n8), .Q(n7) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n5) );
  AO222X1 U12 ( .IN1(N65), .IN2(net20864), .IN3(net20874), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n5), .Q(product2[50]) );
  INVX0 U3 ( .INP(n3), .ZN(n4) );
  INVX0 U4 ( .INP(product_shift[35]), .ZN(n3) );
  NBUFFX2 U55 ( .INP(n7), .Z(net20874) );
  NBUFFX2 U57 ( .INP(n6), .Z(net20864) );
  NBUFFX2 U60 ( .INP(n5), .Z(net20886) );
  NBUFFX2 U61 ( .INP(n5), .Z(net20888) );
  INVX0 U62 ( .INP(product_shift[0]), .ZN(n8) );
  NOR2X0 U63 ( .IN1(n8), .IN2(product_shift[1]), .QN(n6) );
  INVX0 U64 ( .INP(combined_b[7]), .ZN(n9) );
  INVX0 U65 ( .INP(n9), .ZN(n10) );
  INVX0 U66 ( .INP(combined_negative_b[8]), .ZN(n11) );
  INVX0 U67 ( .INP(n11), .ZN(n12) );
  INVX0 U68 ( .INP(product_shift[34]), .ZN(n13) );
  INVX0 U69 ( .INP(n13), .ZN(n14) );
  INVX0 U70 ( .INP(combined_b[6]), .ZN(n15) );
  INVX0 U71 ( .INP(n15), .ZN(n16) );
  INVX0 U72 ( .INP(combined_negative_b[7]), .ZN(n17) );
  INVX0 U73 ( .INP(n17), .ZN(n18) );
  INVX0 U74 ( .INP(product_shift[33]), .ZN(n19) );
  INVX0 U75 ( .INP(n19), .ZN(n20) );
  INVX0 U76 ( .INP(combined_b[5]), .ZN(n21) );
  INVX0 U77 ( .INP(n21), .ZN(n22) );
  INVX0 U78 ( .INP(combined_negative_b[6]), .ZN(n23) );
  INVX0 U79 ( .INP(n23), .ZN(n24) );
  INVX0 U80 ( .INP(product_shift[32]), .ZN(n25) );
  INVX0 U81 ( .INP(n25), .ZN(n26) );
  INVX0 U82 ( .INP(combined_b[4]), .ZN(n27) );
  INVX0 U83 ( .INP(n27), .ZN(n28) );
  INVX0 U84 ( .INP(combined_negative_b[5]), .ZN(n29) );
  INVX0 U85 ( .INP(n29), .ZN(n30) );
  INVX0 U86 ( .INP(product_shift[31]), .ZN(n31) );
  INVX0 U87 ( .INP(n31), .ZN(n32) );
  INVX0 U88 ( .INP(combined_b[3]), .ZN(n33) );
  INVX0 U89 ( .INP(n33), .ZN(n34) );
  INVX0 U90 ( .INP(combined_negative_b[4]), .ZN(n35) );
  INVX0 U91 ( .INP(n35), .ZN(n36) );
  INVX0 U92 ( .INP(product_shift[30]), .ZN(n37) );
  INVX0 U93 ( .INP(n37), .ZN(n38) );
  INVX0 U94 ( .INP(combined_b[2]), .ZN(n39) );
  INVX0 U95 ( .INP(n39), .ZN(n40) );
  INVX0 U96 ( .INP(combined_negative_b[3]), .ZN(n41) );
  INVX0 U97 ( .INP(n41), .ZN(n42) );
  INVX0 U98 ( .INP(product_shift[29]), .ZN(n43) );
  INVX0 U99 ( .INP(n43), .ZN(n44) );
  INVX0 U100 ( .INP(combined_negative_b[2]), .ZN(n45) );
  INVX0 U101 ( .INP(n45), .ZN(n46) );
  INVX0 U102 ( .INP(product_shift[28]), .ZN(n47) );
  INVX0 U103 ( .INP(n47), .ZN(n48) );
  INVX0 U104 ( .INP(combined_negative_b[1]), .ZN(n49) );
  INVX0 U105 ( .INP(n49), .ZN(n50) );
  NBUFFX2 U106 ( .INP(n55), .Z(n56) );
  NBUFFX2 U107 ( .INP(n55), .Z(n57) );
  NBUFFX2 U108 ( .INP(n55), .Z(n58) );
  NBUFFX2 U109 ( .INP(n55), .Z(n59) );
  NBUFFX2 U110 ( .INP(n55), .Z(n60) );
  NBUFFX2 U111 ( .INP(n55), .Z(n61) );
  NBUFFX2 U112 ( .INP(n55), .Z(n62) );
  NBUFFX2 U113 ( .INP(n55), .Z(n63) );
  NBUFFX2 U114 ( .INP(n55), .Z(n65) );
  NBUFFX2 U115 ( .INP(n55), .Z(n66) );
  NBUFFX2 U116 ( .INP(n55), .Z(n67) );
  NBUFFX2 U117 ( .INP(n55), .Z(n64) );
  NBUFFX2 U118 ( .INP(n6), .Z(net20870) );
  NBUFFX2 U119 ( .INP(n6), .Z(net20868) );
  NBUFFX2 U120 ( .INP(n6), .Z(net20866) );
  NBUFFX2 U121 ( .INP(n7), .Z(net20876) );
  NBUFFX2 U122 ( .INP(reset), .Z(n55) );
  INVX0 U124 ( .INP(product_shift[27]), .ZN(n51) );
  INVX0 U125 ( .INP(n51), .ZN(n52) );
  INVX0 U126 ( .INP(product_shift[26]), .ZN(n53) );
  INVX0 U127 ( .INP(n53), .ZN(n54) );
endmodule


module booth6_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n24), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1 ( .IN1(A[30]), .IN2(B[30]), .IN3(carry[30]), .Q(SUM[30]) );
  XOR2X1 U2 ( .IN1(A[31]), .IN2(B[31]), .Q(n17) );
  XOR3X1 U3 ( .IN1(A[42]), .IN2(B[42]), .IN3(carry[42]), .Q(SUM[42]) );
  NAND2X0 U4 ( .IN1(A[42]), .IN2(B[42]), .QN(n1) );
  NAND2X0 U5 ( .IN1(A[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X0 U6 ( .IN1(B[42]), .IN2(carry[42]), .QN(n3) );
  NAND3X0 U7 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[43]) );
  XOR2X1 U8 ( .IN1(A[43]), .IN2(B[43]), .Q(n4) );
  XOR2X1 U9 ( .IN1(n4), .IN2(carry[43]), .Q(SUM[43]) );
  NAND2X0 U10 ( .IN1(A[43]), .IN2(B[43]), .QN(n5) );
  NAND2X0 U11 ( .IN1(A[43]), .IN2(carry[43]), .QN(n6) );
  NAND2X0 U12 ( .IN1(B[43]), .IN2(carry[43]), .QN(n7) );
  NAND3X0 U13 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[44]) );
  XOR3X1 U14 ( .IN1(carry[34]), .IN2(B[34]), .IN3(A[34]), .Q(SUM[34]) );
  NAND2X0 U15 ( .IN1(A[34]), .IN2(carry[34]), .QN(n8) );
  NAND2X0 U16 ( .IN1(B[34]), .IN2(carry[34]), .QN(n9) );
  NAND2X0 U17 ( .IN1(B[34]), .IN2(A[34]), .QN(n10) );
  NAND3X0 U18 ( .IN1(n8), .IN2(n10), .IN3(n9), .QN(carry[35]) );
  XOR3X1 U19 ( .IN1(carry[41]), .IN2(B[41]), .IN3(A[41]), .Q(SUM[41]) );
  NAND2X0 U20 ( .IN1(A[41]), .IN2(carry[41]), .QN(n11) );
  NAND2X0 U21 ( .IN1(B[41]), .IN2(carry[41]), .QN(n12) );
  NAND2X0 U22 ( .IN1(B[41]), .IN2(A[41]), .QN(n13) );
  NAND3X0 U23 ( .IN1(n11), .IN2(n13), .IN3(n12), .QN(carry[42]) );
  NAND2X0 U24 ( .IN1(A[30]), .IN2(B[30]), .QN(n14) );
  NAND2X0 U25 ( .IN1(A[30]), .IN2(carry[30]), .QN(n15) );
  NAND2X0 U26 ( .IN1(B[30]), .IN2(carry[30]), .QN(n16) );
  NAND3X0 U27 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[31]) );
  XOR2X1 U28 ( .IN1(n17), .IN2(carry[31]), .Q(SUM[31]) );
  NAND2X0 U29 ( .IN1(A[31]), .IN2(B[31]), .QN(n18) );
  NAND2X0 U30 ( .IN1(A[31]), .IN2(carry[31]), .QN(n19) );
  NAND2X0 U31 ( .IN1(B[31]), .IN2(carry[31]), .QN(n20) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[32]) );
  XOR3X1 U33 ( .IN1(carry[35]), .IN2(A[35]), .IN3(B[35]), .Q(SUM[35]) );
  NAND2X0 U34 ( .IN1(B[35]), .IN2(carry[35]), .QN(n21) );
  NAND2X0 U35 ( .IN1(A[35]), .IN2(carry[35]), .QN(n22) );
  NAND2X0 U36 ( .IN1(A[35]), .IN2(B[35]), .QN(n23) );
  NAND3X0 U37 ( .IN1(n21), .IN2(n23), .IN3(n22), .QN(carry[36]) );
  AND2X1 U38 ( .IN1(A[26]), .IN2(B[26]), .Q(n24) );
  XOR2X1 U39 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_10_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X1 U1 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X1 U2 ( .IN1(A[46]), .IN2(carry[46]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[46]), .IN2(carry[46]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[46]), .IN2(A[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[47]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  XOR3X1 U7 ( .IN1(B[35]), .IN2(A[35]), .IN3(carry[35]), .Q(SUM[35]) );
  NAND2X1 U8 ( .IN1(carry[35]), .IN2(B[35]), .QN(n4) );
  NAND2X1 U9 ( .IN1(A[35]), .IN2(B[35]), .QN(n5) );
  NAND2X0 U10 ( .IN1(A[35]), .IN2(carry[35]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[36]) );
  INVX0 U12 ( .INP(carry[48]), .ZN(n7) );
  INVX0 U13 ( .INP(n7), .ZN(n8) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n9) );
  XOR3X1 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X1 U16 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  AND2X1 U17 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  NAND2X0 U18 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U22 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U24 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U28 ( .IN1(n16), .IN2(n15), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U34 ( .IN1(n20), .IN2(n8), .Q(SUM[48]) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U40 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U41 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_10 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N24, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[10] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n76), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n76), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n75), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n72), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n71), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n71), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n70), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n70), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n69), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n69), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n11), .CLK(clk), .RSTB(n69), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n17), .CLK(clk), .RSTB(n69), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n23), .CLK(clk), .RSTB(n69), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n29), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n35), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n41), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n45), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n49), .CLK(clk), .RSTB(n68), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n68), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n68), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n67), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n67), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n67), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n66), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n65), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n65), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n65), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n65), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n65), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n65), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n65), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n65), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n65), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n65), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n61), .IN3(N75), .IN4(n57), .IN5(
        product_shift[9]), .IN6(n55), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n61), .IN3(N74), .IN4(n57), .IN5(
        product_shift[8]), .IN6(n78), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n61), .IN3(N73), .IN4(n57), .IN5(
        product_shift[7]), .IN6(n78), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n61), .IN3(N72), .IN4(n57), .IN5(
        product_shift[6]), .IN6(n56), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n61), .IN3(N71), .IN4(n57), .IN5(
        product_shift[5]), .IN6(n78), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n61), .IN3(n57), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n56), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n61), .IN3(N70), .IN4(n57), .IN5(
        product_shift[4]), .IN6(n55), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n61), .IN3(N115), .IN4(n57), .IN5(
        product_shift[49]), .IN6(n78), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n61), .IN3(N114), .IN4(n57), .IN5(
        product_shift[48]), .IN6(n78), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n61), .IN3(N113), .IN4(n57), .IN5(
        product_shift[47]), .IN6(n78), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n61), .IN3(N112), .IN4(n57), .IN5(
        product_shift[46]), .IN6(n78), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n61), .IN3(N111), .IN4(n57), .IN5(
        product_shift[45]), .IN6(n78), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n62), .IN3(N110), .IN4(n58), .IN5(
        product_shift[44]), .IN6(n56), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n62), .IN3(N109), .IN4(n58), .IN5(
        product_shift[43]), .IN6(n56), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n62), .IN3(N108), .IN4(n58), .IN5(
        product_shift[42]), .IN6(n56), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n62), .IN3(N107), .IN4(n58), .IN5(
        product_shift[41]), .IN6(n56), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n62), .IN3(N106), .IN4(n58), .IN5(
        product_shift[40]), .IN6(n56), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n62), .IN3(N69), .IN4(n58), .IN5(
        product_shift[3]), .IN6(n56), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n62), .IN3(N105), .IN4(n58), .IN5(
        product_shift[39]), .IN6(n56), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n62), .IN3(N104), .IN4(n58), .IN5(
        product_shift[38]), .IN6(n56), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n62), .IN3(N103), .IN4(n58), .IN5(
        product_shift[37]), .IN6(n56), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n62), .IN3(N102), .IN4(n58), .IN5(
        product_shift[36]), .IN6(n56), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n62), .IN3(N101), .IN4(n58), .IN5(n4), .IN6(
        n56), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n62), .IN3(N100), .IN4(n58), .IN5(n13), .IN6(
        n56), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n63), .IN3(N99), .IN4(n59), .IN5(n19), .IN6(
        n56), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n63), .IN3(N98), .IN4(n59), .IN5(n25), .IN6(
        n55), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n63), .IN3(N97), .IN4(n59), .IN5(n31), .IN6(
        n78), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n63), .IN3(N96), .IN4(n59), .IN5(n37), .IN6(
        n78), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n63), .IN3(N68), .IN4(n59), .IN5(
        product_shift[2]), .IN6(n78), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n63), .IN3(N95), .IN4(n59), .IN5(n43), .IN6(
        n78), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n63), .IN3(N94), .IN4(n59), .IN5(n47), .IN6(
        n78), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n63), .IN3(N93), .IN4(n59), .IN5(n51), .IN6(
        n78), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n63), .IN3(N92), .IN4(n59), .IN5(n53), .IN6(
        n78), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n63), .IN3(N91), .IN4(n59), .IN5(
        product_shift[25]), .IN6(n78), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n63), .IN3(N90), .IN4(n59), .IN5(
        product_shift[24]), .IN6(n78), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n63), .IN3(N89), .IN4(n59), .IN5(
        product_shift[23]), .IN6(n78), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n64), .IN3(N88), .IN4(n60), .IN5(
        product_shift[22]), .IN6(n56), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n64), .IN3(N87), .IN4(n60), .IN5(
        product_shift[21]), .IN6(n55), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n64), .IN3(N86), .IN4(n60), .IN5(
        product_shift[20]), .IN6(n55), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n64), .IN3(N67), .IN4(n60), .IN5(n55), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n64), .IN3(N85), .IN4(n60), .IN5(
        product_shift[19]), .IN6(n55), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n64), .IN3(N84), .IN4(n60), .IN5(
        product_shift[18]), .IN6(n55), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n64), .IN3(N83), .IN4(n60), .IN5(
        product_shift[17]), .IN6(n55), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n64), .IN3(N82), .IN4(n60), .IN5(
        product_shift[16]), .IN6(n55), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n64), .IN3(N81), .IN4(n60), .IN5(
        product_shift[15]), .IN6(n55), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n64), .IN3(N80), .IN4(n60), .IN5(
        product_shift[14]), .IN6(n55), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n64), .IN3(N79), .IN4(n60), .IN5(
        product_shift[13]), .IN6(n55), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n64), .IN3(N78), .IN4(n60), .IN5(
        product_shift[12]), .IN6(n55), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n64), .IN3(N77), .IN4(n60), .IN5(
        product_shift[11]), .IN6(n55), .Q(product2[11]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n78) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n77), .Q(n79) );
  booth6_10_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], 
        n4, n13, n19, n25, n31, n37, n43, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_negative_b[24:9], n11, n17, n23, n29, n35, n41, n45, n49, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        SYNOPSYS_UNCONNECTED__0, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_10_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:36], 
        n4, n13, n19, n25, n31, n37, n43, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, SYNOPSYS_UNCONNECTED__2, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(n10), .ZN(n11) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U56 ( .INP(product_shift[35]), .ZN(n3) );
  INVX0 U57 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U60 ( .INP(n5), .ZN(n9) );
  INVX0 U61 ( .INP(combined_negative_b[8]), .ZN(n10) );
  INVX0 U62 ( .INP(product_shift[34]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(combined_negative_b[7]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(product_shift[33]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(combined_negative_b[6]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(product_shift[32]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(combined_negative_b[5]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(product_shift[31]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(combined_negative_b[4]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(product_shift[30]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(combined_negative_b[3]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(product_shift[29]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_negative_b[2]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  INVX0 U96 ( .INP(product_shift[28]), .ZN(n46) );
  INVX0 U97 ( .INP(n46), .ZN(n47) );
  INVX0 U98 ( .INP(combined_negative_b[1]), .ZN(n48) );
  INVX0 U99 ( .INP(n48), .ZN(n49) );
  NBUFFX2 U100 ( .INP(n54), .Z(n65) );
  NBUFFX2 U101 ( .INP(n54), .Z(n66) );
  NBUFFX2 U102 ( .INP(n54), .Z(n67) );
  NBUFFX2 U103 ( .INP(n54), .Z(n68) );
  NBUFFX2 U104 ( .INP(n54), .Z(n69) );
  NBUFFX2 U105 ( .INP(n54), .Z(n70) );
  NBUFFX2 U106 ( .INP(n54), .Z(n71) );
  NBUFFX2 U107 ( .INP(n54), .Z(n72) );
  NBUFFX2 U108 ( .INP(n54), .Z(n74) );
  NBUFFX2 U109 ( .INP(n54), .Z(n75) );
  NBUFFX2 U110 ( .INP(n54), .Z(n76) );
  NBUFFX2 U111 ( .INP(n54), .Z(n73) );
  NBUFFX2 U112 ( .INP(n80), .Z(n64) );
  NBUFFX2 U113 ( .INP(n80), .Z(n63) );
  NBUFFX2 U114 ( .INP(n80), .Z(n62) );
  NBUFFX2 U115 ( .INP(n80), .Z(n61) );
  NBUFFX2 U116 ( .INP(n78), .Z(n55) );
  NBUFFX2 U117 ( .INP(n78), .Z(n56) );
  NBUFFX2 U118 ( .INP(n79), .Z(n60) );
  NBUFFX2 U119 ( .INP(n79), .Z(n59) );
  NBUFFX2 U120 ( .INP(n79), .Z(n58) );
  NBUFFX2 U121 ( .INP(n79), .Z(n57) );
  NBUFFX2 U122 ( .INP(reset), .Z(n54) );
  NOR2X0 U123 ( .IN1(n77), .IN2(product_shift[1]), .QN(n80) );
  INVX0 U124 ( .INP(product_shift[0]), .ZN(n77) );
  INVX0 U126 ( .INP(product_shift[27]), .ZN(n50) );
  INVX0 U127 ( .INP(n50), .ZN(n51) );
  INVX0 U128 ( .INP(product_shift[26]), .ZN(n52) );
  INVX0 U129 ( .INP(n52), .ZN(n53) );
endmodule


module booth6_9_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n41), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX2 U1_35 ( .A(carry[35]), .B(B[35]), .CI(A[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[47]), .IN2(B[47]), .IN3(A[47]), .Q(SUM[47]) );
  NAND2X1 U2 ( .IN1(A[47]), .IN2(carry[47]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[47]), .IN2(carry[47]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[47]), .IN2(A[47]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[48]) );
  XOR3X1 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  XOR3X1 U7 ( .IN1(A[40]), .IN2(B[40]), .IN3(n12), .Q(SUM[40]) );
  XOR3X1 U8 ( .IN1(A[43]), .IN2(B[43]), .IN3(n11), .Q(SUM[43]) );
  NAND2X0 U9 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U10 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U11 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U12 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U13 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U14 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U15 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U16 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U17 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U18 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  DELLN2X2 U19 ( .INP(carry[43]), .Z(n11) );
  DELLN2X2 U20 ( .INP(carry[40]), .Z(n12) );
  XOR3X1 U21 ( .IN1(carry[39]), .IN2(B[39]), .IN3(A[39]), .Q(SUM[39]) );
  NAND2X0 U22 ( .IN1(A[39]), .IN2(carry[39]), .QN(n13) );
  NAND2X0 U23 ( .IN1(B[39]), .IN2(carry[39]), .QN(n14) );
  NAND2X0 U24 ( .IN1(B[39]), .IN2(A[39]), .QN(n15) );
  NAND3X0 U25 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[40]) );
  DELLN2X2 U26 ( .INP(carry[46]), .Z(n16) );
  DELLN2X2 U27 ( .INP(carry[44]), .Z(n17) );
  XOR3X1 U28 ( .IN1(A[45]), .IN2(B[45]), .IN3(n19), .Q(SUM[45]) );
  DELLN2X2 U29 ( .INP(carry[41]), .Z(n18) );
  DELLN2X2 U30 ( .INP(carry[45]), .Z(n19) );
  NAND2X0 U31 ( .IN1(A[45]), .IN2(B[45]), .QN(n20) );
  NAND2X0 U32 ( .IN1(A[45]), .IN2(carry[45]), .QN(n21) );
  NAND2X0 U33 ( .IN1(B[45]), .IN2(carry[45]), .QN(n22) );
  NAND3X0 U34 ( .IN1(n21), .IN2(n22), .IN3(n20), .QN(carry[46]) );
  XOR2X1 U35 ( .IN1(A[46]), .IN2(B[46]), .Q(n23) );
  XOR2X1 U36 ( .IN1(n23), .IN2(n16), .Q(SUM[46]) );
  NAND2X0 U37 ( .IN1(A[46]), .IN2(B[46]), .QN(n24) );
  NAND2X0 U38 ( .IN1(A[46]), .IN2(carry[46]), .QN(n25) );
  NAND2X0 U39 ( .IN1(B[46]), .IN2(carry[46]), .QN(n26) );
  NAND3X0 U40 ( .IN1(n24), .IN2(n25), .IN3(n26), .QN(carry[47]) );
  NAND2X0 U41 ( .IN1(A[43]), .IN2(B[43]), .QN(n27) );
  NAND2X0 U42 ( .IN1(A[43]), .IN2(carry[43]), .QN(n28) );
  NAND2X0 U43 ( .IN1(B[43]), .IN2(carry[43]), .QN(n29) );
  NAND3X0 U44 ( .IN1(n28), .IN2(n29), .IN3(n27), .QN(carry[44]) );
  XOR2X1 U45 ( .IN1(A[44]), .IN2(B[44]), .Q(n30) );
  XOR2X1 U46 ( .IN1(n30), .IN2(n17), .Q(SUM[44]) );
  NAND2X0 U47 ( .IN1(A[44]), .IN2(B[44]), .QN(n31) );
  NAND2X0 U48 ( .IN1(A[44]), .IN2(carry[44]), .QN(n32) );
  NAND2X0 U49 ( .IN1(B[44]), .IN2(carry[44]), .QN(n33) );
  NAND3X0 U50 ( .IN1(n32), .IN2(n33), .IN3(n31), .QN(carry[45]) );
  NAND2X0 U51 ( .IN1(A[40]), .IN2(B[40]), .QN(n34) );
  NAND2X0 U52 ( .IN1(A[40]), .IN2(carry[40]), .QN(n35) );
  NAND2X0 U53 ( .IN1(B[40]), .IN2(carry[40]), .QN(n36) );
  NAND3X0 U54 ( .IN1(n35), .IN2(n36), .IN3(n34), .QN(carry[41]) );
  XOR2X1 U55 ( .IN1(A[41]), .IN2(B[41]), .Q(n37) );
  XOR2X1 U56 ( .IN1(n37), .IN2(n18), .Q(SUM[41]) );
  NAND2X0 U57 ( .IN1(A[41]), .IN2(B[41]), .QN(n38) );
  NAND2X0 U58 ( .IN1(A[41]), .IN2(carry[41]), .QN(n39) );
  NAND2X0 U59 ( .IN1(B[41]), .IN2(carry[41]), .QN(n40) );
  NAND3X0 U60 ( .IN1(n38), .IN2(n39), .IN3(n40), .QN(carry[42]) );
  AND2X1 U61 ( .IN1(A[26]), .IN2(B[26]), .Q(n41) );
  XOR2X1 U62 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_9_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n8), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  XOR3X1 U7 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U8 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  INVX0 U12 ( .INP(A[34]), .ZN(n7) );
  INVX0 U13 ( .INP(n7), .ZN(n8) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n9) );
  XOR3X1 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X1 U16 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  AND2X1 U17 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  NAND2X0 U18 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U22 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U24 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n17), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U34 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U40 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U41 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_9 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N23, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N74, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[9] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n74), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n74), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n43), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n65), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n63), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n63), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n63), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n63), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n63), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n63), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n63), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n63), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n63), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n63), .Q(add_r2[0])
         );
  AO222X1 U8 ( .IN1(N23), .IN2(n58), .IN3(N74), .IN4(n53), .IN5(
        product_shift[8]), .IN6(n52), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n58), .IN3(N73), .IN4(n53), .IN5(
        product_shift[7]), .IN6(n52), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n58), .IN3(N72), .IN4(n53), .IN5(
        product_shift[6]), .IN6(n52), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n58), .IN3(N71), .IN4(n53), .IN5(
        product_shift[5]), .IN6(n52), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(n58), .IN2(N65), .IN3(n53), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n52), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n58), .IN3(N70), .IN4(n53), .IN5(
        product_shift[4]), .IN6(n52), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n58), .IN3(N115), .IN4(n53), .IN5(
        product_shift[49]), .IN6(n52), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n58), .IN3(N114), .IN4(n53), .IN5(
        product_shift[48]), .IN6(n52), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n58), .IN3(N113), .IN4(n53), .IN5(
        product_shift[47]), .IN6(n52), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n58), .IN3(N112), .IN4(n53), .IN5(
        product_shift[46]), .IN6(n52), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n58), .IN3(N111), .IN4(n53), .IN5(
        product_shift[45]), .IN6(n52), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n59), .IN3(N110), .IN4(n54), .IN5(
        product_shift[44]), .IN6(n51), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n59), .IN3(N109), .IN4(n54), .IN5(
        product_shift[43]), .IN6(n51), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n59), .IN3(N108), .IN4(n54), .IN5(
        product_shift[42]), .IN6(n51), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n59), .IN3(N107), .IN4(n54), .IN5(
        product_shift[41]), .IN6(n51), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n59), .IN3(N106), .IN4(n54), .IN5(
        product_shift[40]), .IN6(n51), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n59), .IN3(N69), .IN4(n54), .IN5(
        product_shift[3]), .IN6(n51), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n59), .IN3(N105), .IN4(n54), .IN5(
        product_shift[39]), .IN6(n51), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n59), .IN3(N104), .IN4(n54), .IN5(
        product_shift[38]), .IN6(n51), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n59), .IN3(N103), .IN4(n54), .IN5(
        product_shift[37]), .IN6(n51), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n59), .IN3(N102), .IN4(n54), .IN5(
        product_shift[36]), .IN6(n51), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n59), .IN3(N101), .IN4(n54), .IN5(
        product_shift[35]), .IN6(n51), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n59), .IN3(N100), .IN4(n54), .IN5(
        product_shift[34]), .IN6(n51), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n60), .IN3(N99), .IN4(n55), .IN5(n11), .IN6(
        n51), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n60), .IN3(N98), .IN4(n55), .IN5(n17), .IN6(
        n50), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n60), .IN3(N97), .IN4(n55), .IN5(n23), .IN6(
        n50), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n60), .IN3(N96), .IN4(n55), .IN5(n29), .IN6(
        n50), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n60), .IN3(N68), .IN4(n55), .IN5(
        product_shift[2]), .IN6(n50), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n60), .IN3(N95), .IN4(n55), .IN5(n35), .IN6(
        n50), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n60), .IN3(N94), .IN4(n55), .IN5(n41), .IN6(
        n50), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n60), .IN3(N93), .IN4(n55), .IN5(n45), .IN6(
        n50), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n60), .IN3(N92), .IN4(n55), .IN5(n47), .IN6(
        n50), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n60), .IN3(N91), .IN4(n55), .IN5(
        product_shift[25]), .IN6(n50), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n60), .IN3(N90), .IN4(n55), .IN5(
        product_shift[24]), .IN6(n50), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n60), .IN3(N89), .IN4(n55), .IN5(
        product_shift[23]), .IN6(n50), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n61), .IN3(N88), .IN4(n56), .IN5(
        product_shift[22]), .IN6(n50), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n61), .IN3(N87), .IN4(n56), .IN5(
        product_shift[21]), .IN6(n49), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n61), .IN3(N86), .IN4(n56), .IN5(
        product_shift[20]), .IN6(n49), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n61), .IN3(N67), .IN4(n56), .IN5(n49), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n61), .IN3(N85), .IN4(n56), .IN5(
        product_shift[19]), .IN6(n49), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n61), .IN3(N84), .IN4(n56), .IN5(
        product_shift[18]), .IN6(n49), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n61), .IN3(N83), .IN4(n56), .IN5(
        product_shift[17]), .IN6(n49), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n61), .IN3(N82), .IN4(n56), .IN5(
        product_shift[16]), .IN6(n49), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n61), .IN3(N81), .IN4(n56), .IN5(
        product_shift[15]), .IN6(n49), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n61), .IN3(N80), .IN4(n56), .IN5(
        product_shift[14]), .IN6(n49), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n61), .IN3(N79), .IN4(n56), .IN5(
        product_shift[13]), .IN6(n49), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n61), .IN3(N78), .IN4(n56), .IN5(
        product_shift[12]), .IN6(n49), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n62), .IN3(N77), .IN4(n57), .IN5(
        product_shift[11]), .IN6(n49), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n62), .IN3(N76), .IN4(n57), .IN5(
        product_shift[10]), .IN6(n50), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n76) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n75), .Q(n77) );
  booth6_9_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n45, n47, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        SYNOPSYS_UNCONNECTED__0, N74, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_9_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n45, n47, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, SYNOPSYS_UNCONNECTED__2, N23, N22, N21, N20, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U7 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_negative_b[1]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  NBUFFX2 U94 ( .INP(n48), .Z(n63) );
  NBUFFX2 U95 ( .INP(n48), .Z(n64) );
  NBUFFX2 U96 ( .INP(n48), .Z(n65) );
  NBUFFX2 U97 ( .INP(n48), .Z(n66) );
  NBUFFX2 U98 ( .INP(n48), .Z(n67) );
  NBUFFX2 U99 ( .INP(n48), .Z(n68) );
  NBUFFX2 U100 ( .INP(n48), .Z(n69) );
  NBUFFX2 U101 ( .INP(n48), .Z(n70) );
  NBUFFX2 U102 ( .INP(n48), .Z(n72) );
  NBUFFX2 U103 ( .INP(n48), .Z(n73) );
  NBUFFX2 U104 ( .INP(n48), .Z(n74) );
  NBUFFX2 U105 ( .INP(n48), .Z(n71) );
  NBUFFX2 U106 ( .INP(n78), .Z(n61) );
  NBUFFX2 U107 ( .INP(n78), .Z(n60) );
  NBUFFX2 U108 ( .INP(n78), .Z(n59) );
  NBUFFX2 U109 ( .INP(n78), .Z(n58) );
  NBUFFX2 U110 ( .INP(n78), .Z(n62) );
  NBUFFX2 U111 ( .INP(n76), .Z(n50) );
  NBUFFX2 U112 ( .INP(n76), .Z(n51) );
  NBUFFX2 U113 ( .INP(n76), .Z(n49) );
  NBUFFX2 U114 ( .INP(n76), .Z(n52) );
  NBUFFX2 U115 ( .INP(n77), .Z(n56) );
  NBUFFX2 U116 ( .INP(n77), .Z(n55) );
  NBUFFX2 U117 ( .INP(n77), .Z(n54) );
  NBUFFX2 U118 ( .INP(n77), .Z(n53) );
  NBUFFX2 U119 ( .INP(n77), .Z(n57) );
  NBUFFX2 U120 ( .INP(reset), .Z(n48) );
  NOR2X0 U121 ( .IN1(n75), .IN2(product_shift[1]), .QN(n78) );
  INVX0 U122 ( .INP(product_shift[0]), .ZN(n75) );
  INVX0 U124 ( .INP(product_shift[27]), .ZN(n44) );
  INVX0 U125 ( .INP(n44), .ZN(n45) );
  INVX0 U126 ( .INP(product_shift[26]), .ZN(n46) );
  INVX0 U127 ( .INP(n46), .ZN(n47) );
endmodule


module booth6_8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[39]), .IN2(B[39]), .IN3(A[39]), .Q(SUM[39]) );
  NAND2X0 U2 ( .IN1(A[39]), .IN2(carry[39]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[39]), .IN2(carry[39]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[39]), .IN2(A[39]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[40]) );
  XNOR2X1 U6 ( .IN1(n31), .IN2(n18), .Q(SUM[47]) );
  XOR3X2 U7 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U9 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U12 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U13 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U15 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U16 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U17 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  XOR3X2 U18 ( .IN1(A[41]), .IN2(B[41]), .IN3(carry[41]), .Q(SUM[41]) );
  NAND2X0 U19 ( .IN1(A[41]), .IN2(B[41]), .QN(n11) );
  NAND2X0 U20 ( .IN1(A[41]), .IN2(carry[41]), .QN(n12) );
  NAND2X0 U21 ( .IN1(B[41]), .IN2(carry[41]), .QN(n13) );
  NAND3X0 U22 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[42]) );
  XOR2X1 U23 ( .IN1(A[42]), .IN2(B[42]), .Q(n14) );
  XOR2X1 U24 ( .IN1(n14), .IN2(carry[42]), .Q(SUM[42]) );
  NAND2X0 U25 ( .IN1(A[42]), .IN2(B[42]), .QN(n15) );
  NAND2X0 U26 ( .IN1(A[42]), .IN2(carry[42]), .QN(n16) );
  NAND2X0 U27 ( .IN1(B[42]), .IN2(carry[42]), .QN(n17) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[43]) );
  INVX0 U29 ( .INP(carry[47]), .ZN(n18) );
  AND2X1 U30 ( .IN1(A[26]), .IN2(B[26]), .Q(n38) );
  XOR3X1 U31 ( .IN1(A[46]), .IN2(B[46]), .IN3(n19), .Q(SUM[46]) );
  DELLN2X2 U32 ( .INP(carry[46]), .Z(n19) );
  DELLN2X2 U33 ( .INP(carry[44]), .Z(n20) );
  XOR3X2 U34 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U35 ( .IN1(A[43]), .IN2(B[43]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[43]), .IN2(carry[43]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[43]), .IN2(carry[43]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n23), .IN3(n21), .QN(carry[44]) );
  XOR2X1 U39 ( .IN1(A[44]), .IN2(B[44]), .Q(n24) );
  XOR2X1 U40 ( .IN1(n24), .IN2(n20), .Q(SUM[44]) );
  NAND2X0 U41 ( .IN1(A[44]), .IN2(B[44]), .QN(n25) );
  NAND2X0 U42 ( .IN1(A[44]), .IN2(carry[44]), .QN(n26) );
  NAND2X0 U43 ( .IN1(B[44]), .IN2(carry[44]), .QN(n27) );
  NAND3X0 U44 ( .IN1(n26), .IN2(n27), .IN3(n25), .QN(carry[45]) );
  NAND2X0 U45 ( .IN1(A[46]), .IN2(B[46]), .QN(n28) );
  NAND2X0 U46 ( .IN1(A[46]), .IN2(carry[46]), .QN(n29) );
  NAND2X0 U47 ( .IN1(B[46]), .IN2(carry[46]), .QN(n30) );
  NAND3X0 U48 ( .IN1(n29), .IN2(n30), .IN3(n28), .QN(carry[47]) );
  XOR2X1 U49 ( .IN1(A[47]), .IN2(B[47]), .Q(n31) );
  NAND2X0 U50 ( .IN1(A[47]), .IN2(B[47]), .QN(n32) );
  NAND2X0 U51 ( .IN1(A[47]), .IN2(carry[47]), .QN(n33) );
  NAND2X0 U52 ( .IN1(B[47]), .IN2(carry[47]), .QN(n34) );
  NAND3X0 U53 ( .IN1(n33), .IN2(n34), .IN3(n32), .QN(carry[48]) );
  XOR3X1 U54 ( .IN1(B[27]), .IN2(n38), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U55 ( .IN1(A[27]), .IN2(B[27]), .QN(n35) );
  NAND2X1 U56 ( .IN1(n38), .IN2(B[27]), .QN(n36) );
  NAND2X0 U57 ( .IN1(n38), .IN2(A[27]), .QN(n37) );
  NAND3X0 U58 ( .IN1(n35), .IN2(n37), .IN3(n36), .QN(carry[28]) );
  XOR2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n10), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  XOR3X1 U1 ( .IN1(carry[40]), .IN2(B[40]), .IN3(A[40]), .Q(SUM[40]) );
  NAND2X0 U2 ( .IN1(A[40]), .IN2(carry[40]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[40]), .IN2(carry[40]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[40]), .IN2(A[40]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[41]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n28), .IN3(A[27]), .Q(SUM[27]) );
  XNOR2X1 U7 ( .IN1(n21), .IN2(n7), .Q(SUM[48]) );
  XOR3X1 U8 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U9 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U11 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U12 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  INVX0 U13 ( .INP(carry[48]), .ZN(n7) );
  DELLN2X2 U14 ( .INP(carry[45]), .Z(n8) );
  INVX0 U15 ( .INP(A[34]), .ZN(n9) );
  INVX0 U16 ( .INP(n9), .ZN(n10) );
  XOR3X1 U17 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X1 U18 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  AND2X1 U19 ( .IN1(A[26]), .IN2(B[26]), .Q(n28) );
  NAND2X0 U20 ( .IN1(n28), .IN2(B[27]), .QN(n26) );
  NAND2X0 U21 ( .IN1(A[44]), .IN2(B[44]), .QN(n11) );
  NAND2X0 U22 ( .IN1(A[44]), .IN2(carry[44]), .QN(n12) );
  NAND2X0 U23 ( .IN1(B[44]), .IN2(carry[44]), .QN(n13) );
  NAND3X0 U24 ( .IN1(n13), .IN2(n12), .IN3(n11), .QN(carry[45]) );
  XOR2X1 U25 ( .IN1(A[45]), .IN2(B[45]), .Q(n14) );
  XOR2X1 U26 ( .IN1(n14), .IN2(n8), .Q(SUM[45]) );
  NAND2X0 U27 ( .IN1(A[45]), .IN2(B[45]), .QN(n15) );
  NAND2X0 U28 ( .IN1(A[45]), .IN2(carry[45]), .QN(n16) );
  NAND2X0 U29 ( .IN1(B[45]), .IN2(carry[45]), .QN(n17) );
  NAND3X0 U30 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[46]) );
  NAND2X0 U31 ( .IN1(A[47]), .IN2(B[47]), .QN(n18) );
  NAND2X0 U32 ( .IN1(A[47]), .IN2(carry[47]), .QN(n19) );
  NAND2X0 U33 ( .IN1(B[47]), .IN2(carry[47]), .QN(n20) );
  NAND3X0 U34 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[48]) );
  XOR2X1 U35 ( .IN1(A[48]), .IN2(B[48]), .Q(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(B[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(A[48]), .IN2(carry[48]), .QN(n23) );
  NAND2X0 U38 ( .IN1(B[48]), .IN2(carry[48]), .QN(n24) );
  NAND3X0 U39 ( .IN1(n23), .IN2(n24), .IN3(n22), .QN(carry[49]) );
  NAND2X0 U40 ( .IN1(A[27]), .IN2(B[27]), .QN(n25) );
  NAND2X0 U41 ( .IN1(n28), .IN2(A[27]), .QN(n27) );
  NAND3X0 U42 ( .IN1(n25), .IN2(n27), .IN3(n26), .QN(carry[28]) );
  XOR2X1 U43 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_8 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N22, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N73,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[8] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n70), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n70), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n66), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n65), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n64), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n63), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n63), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n62), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n62), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n62), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n61), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n61), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n59), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n59), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n59), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n59), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n59), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n59), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n59), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n59), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n59), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n59), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n54), .IN3(N75), .IN4(n49), .IN5(
        product_shift[9]), .IN6(n72), .Q(product2[9]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n54), .IN3(N73), .IN4(n49), .IN5(
        product_shift[7]), .IN6(n48), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n54), .IN3(N72), .IN4(n49), .IN5(
        product_shift[6]), .IN6(n48), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n54), .IN3(N71), .IN4(n49), .IN5(
        product_shift[5]), .IN6(n48), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n54), .IN3(n49), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n54), .IN3(N70), .IN4(n49), .IN5(
        product_shift[4]), .IN6(n48), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n54), .IN3(N115), .IN4(n49), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n54), .IN3(N114), .IN4(n49), .IN5(
        product_shift[48]), .IN6(n48), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n54), .IN3(N113), .IN4(n49), .IN5(
        product_shift[47]), .IN6(n48), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n54), .IN3(N112), .IN4(n49), .IN5(
        product_shift[46]), .IN6(n48), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n54), .IN3(N111), .IN4(n49), .IN5(
        product_shift[45]), .IN6(n48), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n55), .IN3(N110), .IN4(n50), .IN5(
        product_shift[44]), .IN6(n47), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n55), .IN3(N109), .IN4(n50), .IN5(
        product_shift[43]), .IN6(n47), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n55), .IN3(N108), .IN4(n50), .IN5(
        product_shift[42]), .IN6(n47), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n55), .IN3(N107), .IN4(n50), .IN5(
        product_shift[41]), .IN6(n47), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n55), .IN3(N106), .IN4(n50), .IN5(
        product_shift[40]), .IN6(n47), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n55), .IN3(N69), .IN4(n50), .IN5(
        product_shift[3]), .IN6(n47), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n55), .IN3(N105), .IN4(n50), .IN5(
        product_shift[39]), .IN6(n47), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n55), .IN3(N104), .IN4(n50), .IN5(
        product_shift[38]), .IN6(n47), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n55), .IN3(N103), .IN4(n50), .IN5(
        product_shift[37]), .IN6(n47), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n55), .IN3(N102), .IN4(n50), .IN5(
        product_shift[36]), .IN6(n47), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n55), .IN3(N101), .IN4(n50), .IN5(
        product_shift[35]), .IN6(n47), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n55), .IN3(N100), .IN4(n50), .IN5(
        product_shift[34]), .IN6(n47), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n56), .IN3(N99), .IN4(n51), .IN5(n11), .IN6(
        n47), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n56), .IN3(N98), .IN4(n51), .IN5(n17), .IN6(
        n48), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n56), .IN3(N97), .IN4(n51), .IN5(n23), .IN6(
        n48), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n56), .IN3(N96), .IN4(n51), .IN5(n29), .IN6(
        n47), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n56), .IN3(N68), .IN4(n51), .IN5(
        product_shift[2]), .IN6(n48), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n56), .IN3(N95), .IN4(n51), .IN5(n35), .IN6(
        n47), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n56), .IN3(N94), .IN4(n51), .IN5(n41), .IN6(
        n48), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n56), .IN3(N93), .IN4(n51), .IN5(n43), .IN6(
        n72), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n56), .IN3(N92), .IN4(n51), .IN5(n45), .IN6(
        n72), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n56), .IN3(N91), .IN4(n51), .IN5(
        product_shift[25]), .IN6(n72), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n56), .IN3(N90), .IN4(n51), .IN5(
        product_shift[24]), .IN6(n72), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n56), .IN3(N89), .IN4(n51), .IN5(
        product_shift[23]), .IN6(n72), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n57), .IN3(N88), .IN4(n52), .IN5(
        product_shift[22]), .IN6(n72), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n57), .IN3(N87), .IN4(n52), .IN5(
        product_shift[21]), .IN6(n47), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n57), .IN3(N86), .IN4(n52), .IN5(
        product_shift[20]), .IN6(n72), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n57), .IN3(N67), .IN4(n52), .IN5(n72), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n57), .IN3(N85), .IN4(n52), .IN5(
        product_shift[19]), .IN6(n72), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n57), .IN3(N84), .IN4(n52), .IN5(
        product_shift[18]), .IN6(n72), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n57), .IN3(N83), .IN4(n52), .IN5(
        product_shift[17]), .IN6(n72), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n57), .IN3(N82), .IN4(n52), .IN5(
        product_shift[16]), .IN6(n72), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n57), .IN3(N81), .IN4(n52), .IN5(
        product_shift[15]), .IN6(n72), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n57), .IN3(N80), .IN4(n52), .IN5(
        product_shift[14]), .IN6(n72), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n57), .IN3(N79), .IN4(n52), .IN5(
        product_shift[13]), .IN6(n72), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n57), .IN3(N78), .IN4(n52), .IN5(
        product_shift[12]), .IN6(n72), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n58), .IN3(N77), .IN4(n53), .IN5(
        product_shift[11]), .IN6(n48), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n58), .IN3(N76), .IN4(n53), .IN5(
        product_shift[10]), .IN6(n48), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n72) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n71), .Q(n73) );
  booth6_8_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, n45, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, 
        combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, SYNOPSYS_UNCONNECTED__0, N73, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_8_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, n45, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, SYNOPSYS_UNCONNECTED__2, N22, N21, N20, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U8 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  NBUFFX2 U92 ( .INP(n46), .Z(n59) );
  NBUFFX2 U93 ( .INP(n46), .Z(n60) );
  NBUFFX2 U94 ( .INP(n46), .Z(n61) );
  NBUFFX2 U95 ( .INP(n46), .Z(n62) );
  NBUFFX2 U96 ( .INP(n46), .Z(n63) );
  NBUFFX2 U97 ( .INP(n46), .Z(n64) );
  NBUFFX2 U98 ( .INP(n46), .Z(n65) );
  NBUFFX2 U99 ( .INP(n46), .Z(n66) );
  NBUFFX2 U100 ( .INP(n46), .Z(n68) );
  NBUFFX2 U101 ( .INP(n46), .Z(n69) );
  NBUFFX2 U102 ( .INP(n46), .Z(n70) );
  NBUFFX2 U103 ( .INP(n46), .Z(n67) );
  NBUFFX2 U104 ( .INP(n74), .Z(n57) );
  NBUFFX2 U105 ( .INP(n74), .Z(n56) );
  NBUFFX2 U106 ( .INP(n74), .Z(n55) );
  NBUFFX2 U107 ( .INP(n74), .Z(n54) );
  NBUFFX2 U108 ( .INP(n74), .Z(n58) );
  NBUFFX2 U109 ( .INP(n72), .Z(n47) );
  NBUFFX2 U110 ( .INP(n72), .Z(n48) );
  NBUFFX2 U111 ( .INP(n73), .Z(n52) );
  NBUFFX2 U112 ( .INP(n73), .Z(n51) );
  NBUFFX2 U113 ( .INP(n73), .Z(n50) );
  NBUFFX2 U114 ( .INP(n73), .Z(n49) );
  NBUFFX2 U115 ( .INP(n73), .Z(n53) );
  NBUFFX2 U116 ( .INP(reset), .Z(n46) );
  NOR2X0 U117 ( .IN1(n71), .IN2(product_shift[1]), .QN(n74) );
  INVX0 U118 ( .INP(product_shift[0]), .ZN(n71) );
  INVX0 U120 ( .INP(product_shift[27]), .ZN(n42) );
  INVX0 U121 ( .INP(n42), .ZN(n43) );
  INVX0 U122 ( .INP(product_shift[26]), .ZN(n44) );
  INVX0 U123 ( .INP(n44), .ZN(n45) );
endmodule


module booth6_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n30), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_36 ( .A(carry[36]), .B(n10), .CI(A[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X2 U1 ( .IN1(A[33]), .IN2(B[33]), .IN3(carry[33]), .Q(SUM[33]) );
  NAND2X0 U2 ( .IN1(A[33]), .IN2(B[33]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[33]), .IN2(carry[33]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[33]), .IN2(carry[33]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[34]) );
  XOR2X2 U6 ( .IN1(A[34]), .IN2(B[34]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[34]), .Q(SUM[34]) );
  NAND2X0 U8 ( .IN1(A[34]), .IN2(B[34]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[34]), .IN2(carry[34]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[34]), .IN2(carry[34]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[35]) );
  XNOR2X1 U12 ( .IN1(n8), .IN2(carry[30]), .Q(SUM[30]) );
  XNOR2X1 U13 ( .IN1(A[30]), .IN2(B[30]), .Q(n8) );
  INVX0 U14 ( .INP(B[36]), .ZN(n9) );
  INVX0 U15 ( .INP(n9), .ZN(n10) );
  XOR3X2 U16 ( .IN1(A[29]), .IN2(B[29]), .IN3(carry[29]), .Q(SUM[29]) );
  NAND2X0 U17 ( .IN1(A[29]), .IN2(B[29]), .QN(n11) );
  NAND2X0 U18 ( .IN1(A[29]), .IN2(carry[29]), .QN(n12) );
  NAND2X0 U19 ( .IN1(B[29]), .IN2(carry[29]), .QN(n13) );
  NAND3X0 U20 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[30]) );
  NAND2X0 U21 ( .IN1(A[30]), .IN2(B[30]), .QN(n14) );
  NAND2X0 U22 ( .IN1(A[30]), .IN2(carry[30]), .QN(n15) );
  NAND2X0 U23 ( .IN1(B[30]), .IN2(carry[30]), .QN(n16) );
  NAND3X0 U24 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[31]) );
  XOR3X1 U25 ( .IN1(carry[28]), .IN2(B[28]), .IN3(A[28]), .Q(SUM[28]) );
  NAND2X0 U26 ( .IN1(A[28]), .IN2(carry[28]), .QN(n17) );
  NAND2X0 U27 ( .IN1(B[28]), .IN2(carry[28]), .QN(n18) );
  NAND2X0 U28 ( .IN1(B[28]), .IN2(A[28]), .QN(n19) );
  NAND3X0 U29 ( .IN1(n17), .IN2(n19), .IN3(n18), .QN(carry[29]) );
  XOR3X1 U30 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  NAND2X1 U31 ( .IN1(A[31]), .IN2(B[31]), .QN(n20) );
  NAND2X1 U32 ( .IN1(A[31]), .IN2(carry[31]), .QN(n21) );
  NAND2X0 U33 ( .IN1(B[31]), .IN2(carry[31]), .QN(n22) );
  NAND3X0 U34 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(carry[32]) );
  XOR2X1 U35 ( .IN1(A[32]), .IN2(B[32]), .Q(n23) );
  XOR2X1 U36 ( .IN1(n23), .IN2(carry[32]), .Q(SUM[32]) );
  NAND2X0 U37 ( .IN1(A[32]), .IN2(B[32]), .QN(n24) );
  NAND2X0 U38 ( .IN1(A[32]), .IN2(carry[32]), .QN(n25) );
  NAND2X0 U39 ( .IN1(B[32]), .IN2(carry[32]), .QN(n26) );
  NAND3X0 U40 ( .IN1(n24), .IN2(n25), .IN3(n26), .QN(carry[33]) );
  XOR3X1 U41 ( .IN1(carry[35]), .IN2(A[35]), .IN3(B[35]), .Q(SUM[35]) );
  NAND2X0 U42 ( .IN1(B[35]), .IN2(carry[35]), .QN(n27) );
  NAND2X0 U43 ( .IN1(A[35]), .IN2(carry[35]), .QN(n28) );
  NAND2X0 U44 ( .IN1(A[35]), .IN2(B[35]), .QN(n29) );
  NAND3X0 U45 ( .IN1(n27), .IN2(n29), .IN3(n28), .QN(carry[36]) );
  AND2X1 U46 ( .IN1(A[26]), .IN2(B[26]), .Q(n30) );
  XOR2X1 U47 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR2X1 U6 ( .IN1(n18), .IN2(carry[48]), .Q(SUM[48]) );
  XOR3X1 U7 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U8 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  DELLN2X2 U12 ( .INP(carry[45]), .Z(n7) );
  XOR3X1 U13 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X1 U14 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X2 U15 ( .IN1(B[27]), .IN2(n25), .IN3(A[27]), .Q(SUM[27]) );
  AND2X1 U16 ( .IN1(A[26]), .IN2(B[26]), .Q(n25) );
  NAND2X0 U17 ( .IN1(n25), .IN2(B[27]), .QN(n23) );
  NAND2X0 U18 ( .IN1(A[44]), .IN2(B[44]), .QN(n8) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(carry[44]), .QN(n9) );
  NAND2X0 U20 ( .IN1(B[44]), .IN2(carry[44]), .QN(n10) );
  NAND3X0 U21 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[45]) );
  XOR2X1 U22 ( .IN1(A[45]), .IN2(B[45]), .Q(n11) );
  XOR2X1 U23 ( .IN1(n11), .IN2(n7), .Q(SUM[45]) );
  NAND2X0 U24 ( .IN1(A[45]), .IN2(B[45]), .QN(n12) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(carry[45]), .QN(n13) );
  NAND2X0 U26 ( .IN1(B[45]), .IN2(carry[45]), .QN(n14) );
  NAND3X0 U27 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U28 ( .IN1(A[47]), .IN2(B[47]), .QN(n15) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(carry[47]), .QN(n16) );
  NAND2X0 U30 ( .IN1(B[47]), .IN2(carry[47]), .QN(n17) );
  NAND3X0 U31 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[48]) );
  XOR2X1 U32 ( .IN1(A[48]), .IN2(B[48]), .Q(n18) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(B[48]), .QN(n19) );
  NAND2X0 U34 ( .IN1(A[48]), .IN2(carry[48]), .QN(n20) );
  NAND2X0 U35 ( .IN1(B[48]), .IN2(carry[48]), .QN(n21) );
  NAND3X0 U36 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[49]) );
  NAND2X0 U37 ( .IN1(A[27]), .IN2(B[27]), .QN(n22) );
  NAND2X0 U38 ( .IN1(n25), .IN2(A[27]), .QN(n24) );
  NAND3X0 U39 ( .IN1(n22), .IN2(n24), .IN3(n23), .QN(carry[28]) );
  XOR2X1 U40 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_7 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N21, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N72, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[7] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n80), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n80), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n80), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n79), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n78), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n77), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n76), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n76), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n75), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n75), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n75), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n75), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n75), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n75), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n74), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n74), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n74), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n74), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n74), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n74), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n73), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n73), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n11), .CLK(clk), .RSTB(n73), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n17), .CLK(clk), .RSTB(n73), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n23), .CLK(clk), .RSTB(n73), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n29), .CLK(clk), .RSTB(n72), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n35), .CLK(clk), .RSTB(n72), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n41), .CLK(clk), .RSTB(n72), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n45), .CLK(clk), .RSTB(n72), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n49), .CLK(clk), .RSTB(n72), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n72), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n72), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n71), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n71), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n71), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n71), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n71), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n70), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n69), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n69), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n69), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n69), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n69), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n69), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n69), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n69), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n69), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n69), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n69), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n69), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n64), .IN3(N75), .IN4(n59), .IN5(
        product_shift[9]), .IN6(n55), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n64), .IN3(N74), .IN4(n59), .IN5(
        product_shift[8]), .IN6(n58), .Q(product2[8]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n64), .IN3(N72), .IN4(n59), .IN5(
        product_shift[6]), .IN6(n58), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n64), .IN3(N71), .IN4(n59), .IN5(
        product_shift[5]), .IN6(n58), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n64), .IN3(n59), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n58), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n64), .IN3(N70), .IN4(n59), .IN5(
        product_shift[4]), .IN6(n58), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n64), .IN3(N115), .IN4(n59), .IN5(
        product_shift[49]), .IN6(n58), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n64), .IN3(N114), .IN4(n59), .IN5(
        product_shift[48]), .IN6(n58), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n64), .IN3(N113), .IN4(n59), .IN5(
        product_shift[47]), .IN6(n58), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n64), .IN3(N112), .IN4(n59), .IN5(
        product_shift[46]), .IN6(n58), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n64), .IN3(N111), .IN4(n59), .IN5(
        product_shift[45]), .IN6(n58), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n65), .IN3(N110), .IN4(n60), .IN5(
        product_shift[44]), .IN6(n57), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n65), .IN3(N109), .IN4(n60), .IN5(
        product_shift[43]), .IN6(n57), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n65), .IN3(N108), .IN4(n60), .IN5(
        product_shift[42]), .IN6(n57), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n65), .IN3(N107), .IN4(n60), .IN5(
        product_shift[41]), .IN6(n57), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n65), .IN3(N106), .IN4(n60), .IN5(
        product_shift[40]), .IN6(n57), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n65), .IN3(N69), .IN4(n60), .IN5(
        product_shift[3]), .IN6(n57), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n65), .IN3(N105), .IN4(n60), .IN5(
        product_shift[39]), .IN6(n57), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n65), .IN3(N104), .IN4(n60), .IN5(
        product_shift[38]), .IN6(n57), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n65), .IN3(N103), .IN4(n60), .IN5(
        product_shift[37]), .IN6(n57), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n65), .IN3(N102), .IN4(n60), .IN5(
        product_shift[36]), .IN6(n57), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n65), .IN3(N101), .IN4(n60), .IN5(n4), .IN6(
        n57), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n65), .IN3(N100), .IN4(n60), .IN5(n13), .IN6(
        n57), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n66), .IN3(N99), .IN4(n61), .IN5(n19), .IN6(
        n57), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n66), .IN3(N98), .IN4(n61), .IN5(n25), .IN6(
        n56), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n66), .IN3(N97), .IN4(n61), .IN5(n31), .IN6(
        n56), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n66), .IN3(N96), .IN4(n61), .IN5(n37), .IN6(
        n56), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n66), .IN3(N68), .IN4(n61), .IN5(
        product_shift[2]), .IN6(n56), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n66), .IN3(N95), .IN4(n61), .IN5(n43), .IN6(
        n56), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n66), .IN3(N94), .IN4(n61), .IN5(n47), .IN6(
        n56), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n66), .IN3(N93), .IN4(n61), .IN5(n51), .IN6(
        n56), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n66), .IN3(N92), .IN4(n61), .IN5(n53), .IN6(
        n56), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n66), .IN3(N91), .IN4(n61), .IN5(
        product_shift[25]), .IN6(n56), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n66), .IN3(N90), .IN4(n61), .IN5(
        product_shift[24]), .IN6(n56), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n66), .IN3(N89), .IN4(n61), .IN5(
        product_shift[23]), .IN6(n56), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n67), .IN3(N88), .IN4(n62), .IN5(
        product_shift[22]), .IN6(n56), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n67), .IN3(N87), .IN4(n62), .IN5(
        product_shift[21]), .IN6(n55), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n67), .IN3(N86), .IN4(n62), .IN5(
        product_shift[20]), .IN6(n55), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n67), .IN3(N67), .IN4(n62), .IN5(n55), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n67), .IN3(N85), .IN4(n62), .IN5(
        product_shift[19]), .IN6(n55), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n67), .IN3(N84), .IN4(n62), .IN5(
        product_shift[18]), .IN6(n55), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n67), .IN3(N83), .IN4(n62), .IN5(
        product_shift[17]), .IN6(n55), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n67), .IN3(N82), .IN4(n62), .IN5(
        product_shift[16]), .IN6(n55), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n67), .IN3(N81), .IN4(n62), .IN5(
        product_shift[15]), .IN6(n55), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n67), .IN3(N80), .IN4(n62), .IN5(
        product_shift[14]), .IN6(n55), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n67), .IN3(N79), .IN4(n62), .IN5(
        product_shift[13]), .IN6(n55), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n67), .IN3(N78), .IN4(n62), .IN5(
        product_shift[12]), .IN6(n55), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n68), .IN3(N77), .IN4(n63), .IN5(
        product_shift[11]), .IN6(n55), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n68), .IN3(N76), .IN4(n63), .IN5(
        product_shift[10]), .IN6(n56), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n82) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n81), .Q(n83) );
  booth6_7_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], n4, 
        n13, n19, n25, n31, n37, n43, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_negative_b[24:9], n11, n17, n23, n29, n35, n41, n45, n49, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, SYNOPSYS_UNCONNECTED__0, N72, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_7_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:36], n4, 
        n13, n19, n25, n31, n37, n43, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, SYNOPSYS_UNCONNECTED__2, N21, N20, 
        N19, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(n3), .ZN(n4) );
  INVX0 U4 ( .INP(n44), .ZN(n45) );
  INVX0 U9 ( .INP(product_shift[35]), .ZN(n3) );
  INVX0 U57 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U60 ( .INP(n5), .ZN(n9) );
  INVX0 U61 ( .INP(combined_negative_b[8]), .ZN(n10) );
  INVX0 U62 ( .INP(n10), .ZN(n11) );
  INVX0 U63 ( .INP(product_shift[34]), .ZN(n12) );
  INVX0 U64 ( .INP(n12), .ZN(n13) );
  INVX0 U65 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U66 ( .INP(n14), .ZN(n15) );
  INVX0 U67 ( .INP(combined_negative_b[7]), .ZN(n16) );
  INVX0 U68 ( .INP(n16), .ZN(n17) );
  INVX0 U69 ( .INP(product_shift[33]), .ZN(n18) );
  INVX0 U70 ( .INP(n18), .ZN(n19) );
  INVX0 U71 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U72 ( .INP(n20), .ZN(n21) );
  INVX0 U73 ( .INP(combined_negative_b[6]), .ZN(n22) );
  INVX0 U74 ( .INP(n22), .ZN(n23) );
  INVX0 U75 ( .INP(product_shift[32]), .ZN(n24) );
  INVX0 U76 ( .INP(n24), .ZN(n25) );
  INVX0 U77 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U78 ( .INP(n26), .ZN(n27) );
  INVX0 U79 ( .INP(combined_negative_b[5]), .ZN(n28) );
  INVX0 U80 ( .INP(n28), .ZN(n29) );
  INVX0 U81 ( .INP(product_shift[31]), .ZN(n30) );
  INVX0 U82 ( .INP(n30), .ZN(n31) );
  INVX0 U83 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U84 ( .INP(n32), .ZN(n33) );
  INVX0 U85 ( .INP(combined_negative_b[4]), .ZN(n34) );
  INVX0 U86 ( .INP(n34), .ZN(n35) );
  INVX0 U87 ( .INP(product_shift[30]), .ZN(n36) );
  INVX0 U88 ( .INP(n36), .ZN(n37) );
  INVX0 U89 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U90 ( .INP(n38), .ZN(n39) );
  INVX0 U91 ( .INP(combined_negative_b[3]), .ZN(n40) );
  INVX0 U92 ( .INP(n40), .ZN(n41) );
  INVX0 U93 ( .INP(product_shift[29]), .ZN(n42) );
  INVX0 U94 ( .INP(n42), .ZN(n43) );
  INVX0 U95 ( .INP(combined_negative_b[2]), .ZN(n44) );
  INVX0 U96 ( .INP(product_shift[28]), .ZN(n46) );
  INVX0 U97 ( .INP(n46), .ZN(n47) );
  INVX0 U98 ( .INP(combined_negative_b[1]), .ZN(n48) );
  INVX0 U99 ( .INP(n48), .ZN(n49) );
  NBUFFX2 U100 ( .INP(n54), .Z(n69) );
  NBUFFX2 U101 ( .INP(n54), .Z(n70) );
  NBUFFX2 U102 ( .INP(n54), .Z(n71) );
  NBUFFX2 U103 ( .INP(n54), .Z(n72) );
  NBUFFX2 U104 ( .INP(n54), .Z(n73) );
  NBUFFX2 U105 ( .INP(n54), .Z(n74) );
  NBUFFX2 U106 ( .INP(n54), .Z(n75) );
  NBUFFX2 U107 ( .INP(n54), .Z(n76) );
  NBUFFX2 U108 ( .INP(n54), .Z(n78) );
  NBUFFX2 U109 ( .INP(n54), .Z(n79) );
  NBUFFX2 U110 ( .INP(n54), .Z(n80) );
  NBUFFX2 U111 ( .INP(n54), .Z(n77) );
  NBUFFX2 U112 ( .INP(n84), .Z(n67) );
  NBUFFX2 U113 ( .INP(n84), .Z(n66) );
  NBUFFX2 U114 ( .INP(n84), .Z(n65) );
  NBUFFX2 U115 ( .INP(n84), .Z(n64) );
  NBUFFX2 U116 ( .INP(n84), .Z(n68) );
  NBUFFX2 U117 ( .INP(n82), .Z(n55) );
  NBUFFX2 U118 ( .INP(n82), .Z(n56) );
  NBUFFX2 U119 ( .INP(n82), .Z(n57) );
  NBUFFX2 U120 ( .INP(n82), .Z(n58) );
  NBUFFX2 U121 ( .INP(n83), .Z(n62) );
  NBUFFX2 U122 ( .INP(n83), .Z(n61) );
  NBUFFX2 U123 ( .INP(n83), .Z(n60) );
  NBUFFX2 U124 ( .INP(n83), .Z(n59) );
  NBUFFX2 U125 ( .INP(n83), .Z(n63) );
  NBUFFX2 U126 ( .INP(reset), .Z(n54) );
  NOR2X0 U127 ( .IN1(n81), .IN2(product_shift[1]), .QN(n84) );
  INVX0 U128 ( .INP(product_shift[0]), .ZN(n81) );
  INVX0 U130 ( .INP(product_shift[27]), .ZN(n50) );
  INVX0 U131 ( .INP(n50), .ZN(n51) );
  INVX0 U132 ( .INP(product_shift[26]), .ZN(n52) );
  INVX0 U133 ( .INP(n52), .ZN(n53) );
endmodule


module booth6_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  XOR3X1 U1 ( .IN1(carry[40]), .IN2(B[40]), .IN3(A[40]), .Q(SUM[40]) );
  NAND2X0 U2 ( .IN1(A[40]), .IN2(carry[40]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[40]), .IN2(carry[40]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[40]), .IN2(A[40]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[41]) );
  XOR3X2 U6 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U7 ( .IN1(A[48]), .IN2(B[48]), .QN(n4) );
  NAND2X0 U8 ( .IN1(A[48]), .IN2(carry[48]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[48]), .IN2(carry[48]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[49]) );
  XOR2X1 U11 ( .IN1(A[49]), .IN2(B[49]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U13 ( .IN1(A[49]), .IN2(B[49]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[49]), .IN2(carry[49]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[49]), .IN2(carry[49]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[50]) );
  XOR3X1 U17 ( .IN1(carry[45]), .IN2(B[45]), .IN3(A[45]), .Q(SUM[45]) );
  NAND2X0 U18 ( .IN1(A[45]), .IN2(carry[45]), .QN(n11) );
  NAND2X0 U19 ( .IN1(B[45]), .IN2(carry[45]), .QN(n12) );
  NAND2X0 U20 ( .IN1(B[45]), .IN2(A[45]), .QN(n13) );
  NAND3X0 U21 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[46]) );
  XOR3X1 U22 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U23 ( .IN1(A[42]), .IN2(carry[42]), .QN(n14) );
  NAND2X0 U24 ( .IN1(B[42]), .IN2(carry[42]), .QN(n15) );
  NAND2X0 U25 ( .IN1(B[42]), .IN2(A[42]), .QN(n16) );
  NAND3X0 U26 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[43]) );
  DELLN2X2 U27 ( .INP(carry[47]), .Z(n17) );
  AND2X1 U28 ( .IN1(A[26]), .IN2(B[26]), .Q(n37) );
  XOR3X1 U29 ( .IN1(A[46]), .IN2(B[46]), .IN3(n18), .Q(SUM[46]) );
  DELLN2X2 U30 ( .INP(carry[46]), .Z(n18) );
  DELLN2X2 U31 ( .INP(carry[44]), .Z(n19) );
  XOR3X2 U32 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U33 ( .IN1(A[43]), .IN2(B[43]), .QN(n20) );
  NAND2X0 U34 ( .IN1(A[43]), .IN2(carry[43]), .QN(n21) );
  NAND2X0 U35 ( .IN1(B[43]), .IN2(carry[43]), .QN(n22) );
  NAND3X0 U36 ( .IN1(n21), .IN2(n22), .IN3(n20), .QN(carry[44]) );
  XOR2X1 U37 ( .IN1(A[44]), .IN2(B[44]), .Q(n23) );
  XOR2X1 U38 ( .IN1(n23), .IN2(n19), .Q(SUM[44]) );
  NAND2X0 U39 ( .IN1(A[44]), .IN2(B[44]), .QN(n24) );
  NAND2X0 U40 ( .IN1(A[44]), .IN2(carry[44]), .QN(n25) );
  NAND2X0 U41 ( .IN1(B[44]), .IN2(carry[44]), .QN(n26) );
  NAND3X0 U42 ( .IN1(n25), .IN2(n26), .IN3(n24), .QN(carry[45]) );
  NAND2X0 U43 ( .IN1(A[46]), .IN2(B[46]), .QN(n27) );
  NAND2X0 U44 ( .IN1(A[46]), .IN2(carry[46]), .QN(n28) );
  NAND2X0 U45 ( .IN1(B[46]), .IN2(carry[46]), .QN(n29) );
  NAND3X0 U46 ( .IN1(n28), .IN2(n29), .IN3(n27), .QN(carry[47]) );
  XOR2X1 U47 ( .IN1(A[47]), .IN2(B[47]), .Q(n30) );
  XOR2X1 U48 ( .IN1(n30), .IN2(n17), .Q(SUM[47]) );
  NAND2X0 U49 ( .IN1(A[47]), .IN2(B[47]), .QN(n31) );
  NAND2X0 U50 ( .IN1(A[47]), .IN2(carry[47]), .QN(n32) );
  NAND2X0 U51 ( .IN1(B[47]), .IN2(carry[47]), .QN(n33) );
  NAND3X0 U52 ( .IN1(n32), .IN2(n33), .IN3(n31), .QN(carry[48]) );
  XOR3X1 U53 ( .IN1(B[27]), .IN2(n37), .IN3(A[27]), .Q(SUM[27]) );
  NAND2X0 U54 ( .IN1(A[27]), .IN2(B[27]), .QN(n34) );
  NAND2X1 U55 ( .IN1(n37), .IN2(B[27]), .QN(n35) );
  NAND2X0 U56 ( .IN1(n37), .IN2(A[27]), .QN(n36) );
  NAND3X0 U57 ( .IN1(n34), .IN2(n36), .IN3(n35), .QN(carry[28]) );
  XOR2X1 U58 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  XOR3X1 U1 ( .IN1(carry[41]), .IN2(B[41]), .IN3(A[41]), .Q(SUM[41]) );
  NAND2X0 U2 ( .IN1(A[41]), .IN2(carry[41]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[41]), .IN2(carry[41]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[41]), .IN2(A[41]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[42]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  XOR3X1 U7 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U8 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U10 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U11 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  DELLN2X2 U12 ( .INP(carry[45]), .Z(n7) );
  INVX0 U13 ( .INP(A[34]), .ZN(n8) );
  INVX0 U14 ( .INP(n8), .ZN(n9) );
  XOR3X2 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X2 U16 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  AND2X1 U17 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  NAND2X0 U18 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U22 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U24 ( .IN1(n13), .IN2(n7), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U28 ( .IN1(n16), .IN2(n15), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U34 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n23), .IN2(n22), .IN3(n21), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U40 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U41 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_6 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N20, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N71, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[6] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n66), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n66), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(combined_negative_b[1]), .CLK(clk), .RSTB(n58), .Q(combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n58), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n57), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n55), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n55), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n55), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n55), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n55), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n55), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n55), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n55), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n55), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n55), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n51), .IN3(N75), .IN4(n49), .IN5(
        product_shift[9]), .IN6(n68), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n51), .IN3(N74), .IN4(n49), .IN5(
        product_shift[8]), .IN6(n48), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n51), .IN3(N73), .IN4(n49), .IN5(
        product_shift[7]), .IN6(n48), .Q(product2[7]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n51), .IN3(N71), .IN4(n49), .IN5(
        product_shift[5]), .IN6(n48), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n51), .IN3(n49), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n51), .IN3(N70), .IN4(n49), .IN5(
        product_shift[4]), .IN6(n48), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n51), .IN3(N115), .IN4(n49), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n51), .IN3(N114), .IN4(n49), .IN5(
        product_shift[48]), .IN6(n48), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n51), .IN3(N113), .IN4(n49), .IN5(
        product_shift[47]), .IN6(n48), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n51), .IN3(N112), .IN4(n49), .IN5(
        product_shift[46]), .IN6(n48), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n51), .IN3(N111), .IN4(n49), .IN5(
        product_shift[45]), .IN6(n48), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n52), .IN3(N110), .IN4(n69), .IN5(
        product_shift[44]), .IN6(n47), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n52), .IN3(N109), .IN4(n69), .IN5(
        product_shift[43]), .IN6(n47), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n52), .IN3(N108), .IN4(n69), .IN5(
        product_shift[42]), .IN6(n47), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n52), .IN3(N107), .IN4(n69), .IN5(
        product_shift[41]), .IN6(n47), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n52), .IN3(N106), .IN4(n69), .IN5(
        product_shift[40]), .IN6(n47), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n52), .IN3(N69), .IN4(n69), .IN5(
        product_shift[3]), .IN6(n47), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n52), .IN3(N105), .IN4(n69), .IN5(
        product_shift[39]), .IN6(n47), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n52), .IN3(N104), .IN4(n69), .IN5(
        product_shift[38]), .IN6(n47), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n52), .IN3(N103), .IN4(n69), .IN5(
        product_shift[37]), .IN6(n47), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n52), .IN3(N102), .IN4(n69), .IN5(
        product_shift[36]), .IN6(n47), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n52), .IN3(N101), .IN4(n69), .IN5(
        product_shift[35]), .IN6(n47), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n52), .IN3(N100), .IN4(n50), .IN5(
        product_shift[34]), .IN6(n47), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n53), .IN3(N99), .IN4(n69), .IN5(n11), .IN6(
        n47), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n53), .IN3(N98), .IN4(n49), .IN5(n17), .IN6(
        n68), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n53), .IN3(N97), .IN4(n50), .IN5(n23), .IN6(
        n68), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n53), .IN3(N96), .IN4(n50), .IN5(n29), .IN6(
        n68), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n53), .IN3(N68), .IN4(n50), .IN5(
        product_shift[2]), .IN6(n68), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n53), .IN3(N95), .IN4(n50), .IN5(n35), .IN6(
        n68), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n53), .IN3(N94), .IN4(n50), .IN5(n41), .IN6(
        n68), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n53), .IN3(N93), .IN4(n50), .IN5(n43), .IN6(
        n48), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n53), .IN3(N92), .IN4(n50), .IN5(n45), .IN6(
        n47), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n53), .IN3(N91), .IN4(n50), .IN5(
        product_shift[25]), .IN6(n48), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n53), .IN3(N90), .IN4(n50), .IN5(
        product_shift[24]), .IN6(n47), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n53), .IN3(N89), .IN4(n50), .IN5(
        product_shift[23]), .IN6(n48), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n53), .IN3(N88), .IN4(n69), .IN5(
        product_shift[22]), .IN6(n48), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n54), .IN3(N87), .IN4(n69), .IN5(
        product_shift[21]), .IN6(n68), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n51), .IN3(N86), .IN4(n69), .IN5(
        product_shift[20]), .IN6(n68), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n54), .IN3(N67), .IN4(n50), .IN5(n68), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n54), .IN3(N85), .IN4(n69), .IN5(
        product_shift[19]), .IN6(n68), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n54), .IN3(N84), .IN4(n69), .IN5(
        product_shift[18]), .IN6(n68), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n54), .IN3(N83), .IN4(n69), .IN5(
        product_shift[17]), .IN6(n68), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n54), .IN3(N82), .IN4(n69), .IN5(
        product_shift[16]), .IN6(n68), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n54), .IN3(N81), .IN4(n69), .IN5(
        product_shift[15]), .IN6(n68), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n54), .IN3(N80), .IN4(n49), .IN5(
        product_shift[14]), .IN6(n68), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n54), .IN3(N79), .IN4(n50), .IN5(
        product_shift[13]), .IN6(n68), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n54), .IN3(N78), .IN4(n49), .IN5(
        product_shift[12]), .IN6(n47), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n54), .IN3(N77), .IN4(n50), .IN5(
        product_shift[11]), .IN6(n48), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n54), .IN3(N76), .IN4(n50), .IN5(
        product_shift[10]), .IN6(n48), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n68) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n67), .Q(n69) );
  booth6_6_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, n45, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, 
        combined_negative_b[1:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        N76, N75, N74, N73, SYNOPSYS_UNCONNECTED__0, N71, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_6_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n43, n45, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, SYNOPSYS_UNCONNECTED__2, N20, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U10 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  NBUFFX2 U92 ( .INP(n46), .Z(n55) );
  NBUFFX2 U93 ( .INP(n46), .Z(n56) );
  NBUFFX2 U94 ( .INP(n46), .Z(n57) );
  NBUFFX2 U95 ( .INP(n46), .Z(n58) );
  NBUFFX2 U96 ( .INP(n46), .Z(n59) );
  NBUFFX2 U97 ( .INP(n46), .Z(n60) );
  NBUFFX2 U98 ( .INP(n46), .Z(n61) );
  NBUFFX2 U99 ( .INP(n46), .Z(n62) );
  NBUFFX2 U100 ( .INP(n46), .Z(n64) );
  NBUFFX2 U101 ( .INP(n46), .Z(n65) );
  NBUFFX2 U102 ( .INP(n46), .Z(n66) );
  NBUFFX2 U103 ( .INP(n46), .Z(n63) );
  NBUFFX2 U104 ( .INP(n70), .Z(n53) );
  NBUFFX2 U105 ( .INP(n70), .Z(n52) );
  NBUFFX2 U106 ( .INP(n70), .Z(n51) );
  NBUFFX2 U107 ( .INP(n70), .Z(n54) );
  NBUFFX2 U108 ( .INP(n68), .Z(n47) );
  NBUFFX2 U109 ( .INP(n68), .Z(n48) );
  NBUFFX2 U110 ( .INP(n69), .Z(n49) );
  NBUFFX2 U111 ( .INP(n69), .Z(n50) );
  NBUFFX2 U112 ( .INP(reset), .Z(n46) );
  NOR2X0 U113 ( .IN1(n67), .IN2(product_shift[1]), .QN(n70) );
  INVX0 U114 ( .INP(product_shift[0]), .ZN(n67) );
  INVX0 U116 ( .INP(product_shift[27]), .ZN(n42) );
  INVX0 U117 ( .INP(n42), .ZN(n43) );
  INVX0 U118 ( .INP(product_shift[26]), .ZN(n44) );
  INVX0 U119 ( .INP(n44), .ZN(n45) );
endmodule


module booth6_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n40), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_33 ( .A(B[33]), .B(A[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  XOR3X2 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U6 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U8 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XNOR2X1 U12 ( .IN1(n22), .IN2(n8), .Q(SUM[47]) );
  INVX0 U13 ( .INP(carry[47]), .ZN(n8) );
  DELLN2X2 U14 ( .INP(carry[42]), .Z(n9) );
  XOR3X1 U15 ( .IN1(A[42]), .IN2(B[42]), .IN3(n9), .Q(SUM[42]) );
  XOR3X1 U16 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  DELLN2X2 U17 ( .INP(carry[41]), .Z(n10) );
  DELLN2X2 U18 ( .INP(carry[43]), .Z(n11) );
  NAND2X0 U19 ( .IN1(A[48]), .IN2(B[48]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[48]), .IN2(carry[48]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[48]), .IN2(carry[48]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n13), .IN2(n14), .IN3(n12), .QN(carry[49]) );
  XOR2X1 U23 ( .IN1(A[49]), .IN2(B[49]), .Q(n15) );
  XOR2X1 U24 ( .IN1(n15), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U25 ( .IN1(A[49]), .IN2(B[49]), .QN(n16) );
  NAND2X0 U26 ( .IN1(A[49]), .IN2(carry[49]), .QN(n17) );
  NAND2X0 U27 ( .IN1(B[49]), .IN2(carry[49]), .QN(n18) );
  NAND3X0 U28 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[50]) );
  XOR3X2 U29 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  NAND2X0 U30 ( .IN1(A[46]), .IN2(B[46]), .QN(n19) );
  NAND2X0 U31 ( .IN1(A[46]), .IN2(carry[46]), .QN(n20) );
  NAND2X0 U32 ( .IN1(B[46]), .IN2(carry[46]), .QN(n21) );
  NAND3X0 U33 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[47]) );
  XOR2X1 U34 ( .IN1(A[47]), .IN2(B[47]), .Q(n22) );
  NAND2X0 U35 ( .IN1(A[47]), .IN2(B[47]), .QN(n23) );
  NAND2X0 U36 ( .IN1(A[47]), .IN2(carry[47]), .QN(n24) );
  NAND2X0 U37 ( .IN1(B[47]), .IN2(carry[47]), .QN(n25) );
  NAND3X0 U38 ( .IN1(n23), .IN2(n24), .IN3(n25), .QN(carry[48]) );
  NAND2X0 U39 ( .IN1(A[42]), .IN2(B[42]), .QN(n26) );
  NAND2X0 U40 ( .IN1(A[42]), .IN2(carry[42]), .QN(n27) );
  NAND2X0 U41 ( .IN1(B[42]), .IN2(carry[42]), .QN(n28) );
  NAND3X0 U42 ( .IN1(n26), .IN2(n27), .IN3(n28), .QN(carry[43]) );
  XOR2X1 U43 ( .IN1(A[43]), .IN2(B[43]), .Q(n29) );
  XOR2X1 U44 ( .IN1(n29), .IN2(n11), .Q(SUM[43]) );
  NAND2X0 U45 ( .IN1(A[43]), .IN2(B[43]), .QN(n30) );
  NAND2X0 U46 ( .IN1(A[43]), .IN2(carry[43]), .QN(n31) );
  NAND2X0 U47 ( .IN1(B[43]), .IN2(carry[43]), .QN(n32) );
  NAND3X0 U48 ( .IN1(n30), .IN2(n31), .IN3(n32), .QN(carry[44]) );
  XOR3X2 U49 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  NAND2X0 U50 ( .IN1(A[40]), .IN2(B[40]), .QN(n33) );
  NAND2X0 U51 ( .IN1(A[40]), .IN2(carry[40]), .QN(n34) );
  NAND2X0 U52 ( .IN1(B[40]), .IN2(carry[40]), .QN(n35) );
  NAND3X0 U53 ( .IN1(n34), .IN2(n35), .IN3(n33), .QN(carry[41]) );
  XOR2X1 U54 ( .IN1(A[41]), .IN2(B[41]), .Q(n36) );
  XOR2X1 U55 ( .IN1(n36), .IN2(n10), .Q(SUM[41]) );
  NAND2X0 U56 ( .IN1(A[41]), .IN2(B[41]), .QN(n37) );
  NAND2X0 U57 ( .IN1(A[41]), .IN2(carry[41]), .QN(n38) );
  NAND2X0 U58 ( .IN1(B[41]), .IN2(carry[41]), .QN(n39) );
  NAND3X0 U59 ( .IN1(n37), .IN2(n38), .IN3(n39), .QN(carry[42]) );
  AND2X1 U60 ( .IN1(A[26]), .IN2(B[26]), .Q(n40) );
  XOR2X1 U61 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(carry[34]), .B(n11), .CI(A[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  XOR3X1 U1 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X1 U2 ( .IN1(A[49]), .IN2(carry[49]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[49]), .IN2(carry[49]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[49]), .IN2(A[49]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[50]) );
  XOR3X1 U6 ( .IN1(B[27]), .IN2(n29), .IN3(A[27]), .Q(SUM[27]) );
  XOR3X1 U7 ( .IN1(A[44]), .IN2(B[44]), .IN3(n7), .Q(SUM[44]) );
  XNOR2X1 U8 ( .IN1(n22), .IN2(n8), .Q(SUM[48]) );
  XOR3X1 U9 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U10 ( .IN1(A[46]), .IN2(carry[46]), .QN(n4) );
  NAND2X0 U11 ( .IN1(B[46]), .IN2(carry[46]), .QN(n5) );
  NAND2X0 U12 ( .IN1(B[46]), .IN2(A[46]), .QN(n6) );
  NAND3X0 U13 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[47]) );
  DELLN2X2 U14 ( .INP(carry[44]), .Z(n7) );
  INVX0 U15 ( .INP(carry[48]), .ZN(n8) );
  DELLN2X2 U16 ( .INP(carry[45]), .Z(n9) );
  INVX0 U17 ( .INP(B[34]), .ZN(n10) );
  INVX0 U18 ( .INP(n10), .ZN(n11) );
  XOR3X2 U19 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  AND2X1 U20 ( .IN1(A[26]), .IN2(B[26]), .Q(n29) );
  NAND2X0 U21 ( .IN1(n29), .IN2(B[27]), .QN(n27) );
  NAND2X0 U22 ( .IN1(A[44]), .IN2(B[44]), .QN(n12) );
  NAND2X0 U23 ( .IN1(A[44]), .IN2(carry[44]), .QN(n13) );
  NAND2X0 U24 ( .IN1(B[44]), .IN2(carry[44]), .QN(n14) );
  NAND3X0 U25 ( .IN1(n14), .IN2(n13), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U26 ( .IN1(A[45]), .IN2(B[45]), .Q(n15) );
  XOR2X1 U27 ( .IN1(n15), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U28 ( .IN1(A[45]), .IN2(B[45]), .QN(n16) );
  NAND2X0 U29 ( .IN1(A[45]), .IN2(carry[45]), .QN(n17) );
  NAND2X0 U30 ( .IN1(B[45]), .IN2(carry[45]), .QN(n18) );
  NAND3X0 U31 ( .IN1(n18), .IN2(n17), .IN3(n16), .QN(carry[46]) );
  NAND2X0 U32 ( .IN1(A[47]), .IN2(B[47]), .QN(n19) );
  NAND2X0 U33 ( .IN1(A[47]), .IN2(carry[47]), .QN(n20) );
  NAND2X0 U34 ( .IN1(B[47]), .IN2(carry[47]), .QN(n21) );
  NAND3X0 U35 ( .IN1(n19), .IN2(n20), .IN3(n21), .QN(carry[48]) );
  XOR2X1 U36 ( .IN1(A[48]), .IN2(B[48]), .Q(n22) );
  NAND2X0 U37 ( .IN1(A[48]), .IN2(B[48]), .QN(n23) );
  NAND2X0 U38 ( .IN1(A[48]), .IN2(carry[48]), .QN(n24) );
  NAND2X0 U39 ( .IN1(B[48]), .IN2(carry[48]), .QN(n25) );
  NAND3X0 U40 ( .IN1(n25), .IN2(n24), .IN3(n23), .QN(carry[49]) );
  NAND2X0 U41 ( .IN1(A[27]), .IN2(B[27]), .QN(n26) );
  NAND2X0 U42 ( .IN1(n29), .IN2(A[27]), .QN(n28) );
  NAND3X0 U43 ( .IN1(n26), .IN2(n28), .IN3(n27), .QN(carry[28]) );
  XOR2X1 U44 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_5 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N19, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N70, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[5] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n66), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n66), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n64), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n63), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n62), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n62), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n61), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n61), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n60), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n60), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n59), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(combined_negative_b[7]), .CLK(clk), .RSTB(n59), .Q(combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n4), .CLK(clk), .RSTB(n59), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n13), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n19), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n25), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n31), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n41), .CLK(clk), .RSTB(n58), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n58), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n58), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n57), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n57), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n57), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n56), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n55), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n55), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n55), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n55), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n55), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n55), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n55), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n55), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n55), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n55), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n55), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n51), .IN3(N75), .IN4(n49), .IN5(
        product_shift[9]), .IN6(n68), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n51), .IN3(N74), .IN4(n49), .IN5(
        product_shift[8]), .IN6(n48), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n51), .IN3(N73), .IN4(n49), .IN5(
        product_shift[7]), .IN6(n48), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n51), .IN3(N72), .IN4(n49), .IN5(
        product_shift[6]), .IN6(n48), .Q(product2[6]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n51), .IN3(n49), .IN4(N116), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n51), .IN3(N70), .IN4(n49), .IN5(
        product_shift[4]), .IN6(n48), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n51), .IN3(N115), .IN4(n49), .IN5(
        product_shift[49]), .IN6(n48), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n51), .IN3(N114), .IN4(n49), .IN5(
        product_shift[48]), .IN6(n48), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n51), .IN3(N113), .IN4(n49), .IN5(
        product_shift[47]), .IN6(n48), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n51), .IN3(N112), .IN4(n49), .IN5(
        product_shift[46]), .IN6(n48), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n51), .IN3(N111), .IN4(n49), .IN5(
        product_shift[45]), .IN6(n48), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n52), .IN3(N110), .IN4(n69), .IN5(
        product_shift[44]), .IN6(n47), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n52), .IN3(N109), .IN4(n69), .IN5(
        product_shift[43]), .IN6(n47), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n52), .IN3(N108), .IN4(n69), .IN5(
        product_shift[42]), .IN6(n47), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n52), .IN3(N107), .IN4(n69), .IN5(
        product_shift[41]), .IN6(n47), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n52), .IN3(N106), .IN4(n69), .IN5(
        product_shift[40]), .IN6(n47), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n52), .IN3(N69), .IN4(n69), .IN5(
        product_shift[3]), .IN6(n47), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n52), .IN3(N105), .IN4(n69), .IN5(
        product_shift[39]), .IN6(n47), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n52), .IN3(N104), .IN4(n69), .IN5(
        product_shift[38]), .IN6(n47), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n52), .IN3(N103), .IN4(n69), .IN5(
        product_shift[37]), .IN6(n47), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n52), .IN3(N102), .IN4(n69), .IN5(
        product_shift[36]), .IN6(n47), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n52), .IN3(N101), .IN4(n69), .IN5(
        product_shift[35]), .IN6(n47), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n52), .IN3(N100), .IN4(n50), .IN5(
        product_shift[34]), .IN6(n47), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n53), .IN3(N99), .IN4(n69), .IN5(n11), .IN6(
        n47), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n53), .IN3(N98), .IN4(n49), .IN5(n17), .IN6(
        n68), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n53), .IN3(N97), .IN4(n50), .IN5(n23), .IN6(
        n68), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n53), .IN3(N96), .IN4(n50), .IN5(n29), .IN6(
        n68), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n53), .IN3(N68), .IN4(n50), .IN5(
        product_shift[2]), .IN6(n68), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n53), .IN3(N95), .IN4(n50), .IN5(n35), .IN6(
        n68), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n53), .IN3(N94), .IN4(n50), .IN5(n39), .IN6(
        n68), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n53), .IN3(N93), .IN4(n50), .IN5(n43), .IN6(
        n48), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n53), .IN3(N92), .IN4(n50), .IN5(n45), .IN6(
        n47), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n53), .IN3(N91), .IN4(n50), .IN5(
        product_shift[25]), .IN6(n48), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n53), .IN3(N90), .IN4(n50), .IN5(
        product_shift[24]), .IN6(n47), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n53), .IN3(N89), .IN4(n50), .IN5(
        product_shift[23]), .IN6(n48), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n53), .IN3(N88), .IN4(n69), .IN5(
        product_shift[22]), .IN6(n48), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n54), .IN3(N87), .IN4(n69), .IN5(
        product_shift[21]), .IN6(n68), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n51), .IN3(N86), .IN4(n69), .IN5(
        product_shift[20]), .IN6(n68), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n54), .IN3(N67), .IN4(n50), .IN5(n68), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n54), .IN3(N85), .IN4(n69), .IN5(
        product_shift[19]), .IN6(n68), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n54), .IN3(N84), .IN4(n69), .IN5(
        product_shift[18]), .IN6(n68), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n54), .IN3(N83), .IN4(n69), .IN5(
        product_shift[17]), .IN6(n68), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n54), .IN3(N82), .IN4(n69), .IN5(
        product_shift[16]), .IN6(n68), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n54), .IN3(N81), .IN4(n69), .IN5(
        product_shift[15]), .IN6(n68), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n54), .IN3(N80), .IN4(n49), .IN5(
        product_shift[14]), .IN6(n68), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n54), .IN3(N79), .IN4(n50), .IN5(
        product_shift[13]), .IN6(n68), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n54), .IN3(N78), .IN4(n49), .IN5(
        product_shift[12]), .IN6(n47), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n54), .IN3(N77), .IN4(n50), .IN5(
        product_shift[11]), .IN6(n48), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n54), .IN3(N76), .IN4(n50), .IN5(
        product_shift[10]), .IN6(n48), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n68) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n67), .Q(n69) );
  booth6_5_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n39, n43, n45, product_shift[25:0]}), .B({
        combined_negative_b[24:7], n4, n13, n19, n25, n31, n41, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, SYNOPSYS_UNCONNECTED__0, N70, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_5_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n39, n43, n45, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n37, combined_b[1:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, SYNOPSYS_UNCONNECTED__2, N19, 
        N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(combined_negative_b[6]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U11 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_negative_b[5]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_negative_b[4]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_negative_b[3]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_negative_b[2]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_b[2]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(product_shift[28]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(combined_negative_b[1]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  NBUFFX2 U92 ( .INP(n46), .Z(n55) );
  NBUFFX2 U93 ( .INP(n46), .Z(n56) );
  NBUFFX2 U94 ( .INP(n46), .Z(n57) );
  NBUFFX2 U95 ( .INP(n46), .Z(n58) );
  NBUFFX2 U96 ( .INP(n46), .Z(n59) );
  NBUFFX2 U97 ( .INP(n46), .Z(n60) );
  NBUFFX2 U98 ( .INP(n46), .Z(n61) );
  NBUFFX2 U99 ( .INP(n46), .Z(n62) );
  NBUFFX2 U100 ( .INP(n46), .Z(n64) );
  NBUFFX2 U101 ( .INP(n46), .Z(n65) );
  NBUFFX2 U102 ( .INP(n46), .Z(n66) );
  NBUFFX2 U103 ( .INP(n46), .Z(n63) );
  NBUFFX2 U104 ( .INP(n70), .Z(n53) );
  NBUFFX2 U105 ( .INP(n70), .Z(n52) );
  NBUFFX2 U106 ( .INP(n70), .Z(n51) );
  NBUFFX2 U107 ( .INP(n70), .Z(n54) );
  NBUFFX2 U108 ( .INP(n68), .Z(n47) );
  NBUFFX2 U109 ( .INP(n68), .Z(n48) );
  NBUFFX2 U110 ( .INP(n69), .Z(n49) );
  NBUFFX2 U111 ( .INP(n69), .Z(n50) );
  NBUFFX2 U112 ( .INP(reset), .Z(n46) );
  NOR2X0 U113 ( .IN1(n67), .IN2(product_shift[1]), .QN(n70) );
  INVX0 U114 ( .INP(product_shift[0]), .ZN(n67) );
  INVX0 U116 ( .INP(product_shift[27]), .ZN(n42) );
  INVX0 U117 ( .INP(n42), .ZN(n43) );
  INVX0 U118 ( .INP(product_shift[26]), .ZN(n44) );
  INVX0 U119 ( .INP(n44), .ZN(n45) );
endmodule


module booth6_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n28), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1 ( .IN1(carry[46]), .IN2(B[46]), .IN3(A[46]), .Q(SUM[46]) );
  NAND2X0 U2 ( .IN1(A[46]), .IN2(carry[46]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[46]), .IN2(carry[46]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[46]), .IN2(A[46]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[47]) );
  XOR3X1 U6 ( .IN1(A[30]), .IN2(B[30]), .IN3(carry[30]), .Q(SUM[30]) );
  XOR2X1 U7 ( .IN1(A[31]), .IN2(B[31]), .Q(n14) );
  XOR3X2 U8 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  NAND2X0 U9 ( .IN1(A[40]), .IN2(B[40]), .QN(n4) );
  NAND2X0 U10 ( .IN1(A[40]), .IN2(carry[40]), .QN(n5) );
  NAND2X0 U11 ( .IN1(B[40]), .IN2(carry[40]), .QN(n6) );
  NAND3X0 U12 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[41]) );
  XOR2X1 U13 ( .IN1(A[41]), .IN2(B[41]), .Q(n7) );
  XOR2X1 U14 ( .IN1(n7), .IN2(carry[41]), .Q(SUM[41]) );
  NAND2X0 U15 ( .IN1(A[41]), .IN2(B[41]), .QN(n8) );
  NAND2X0 U16 ( .IN1(A[41]), .IN2(carry[41]), .QN(n9) );
  NAND2X0 U17 ( .IN1(B[41]), .IN2(carry[41]), .QN(n10) );
  NAND3X0 U18 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[42]) );
  NAND2X0 U19 ( .IN1(A[30]), .IN2(B[30]), .QN(n11) );
  NAND2X0 U20 ( .IN1(A[30]), .IN2(carry[30]), .QN(n12) );
  NAND2X0 U21 ( .IN1(B[30]), .IN2(carry[30]), .QN(n13) );
  NAND3X0 U22 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[31]) );
  XOR2X1 U23 ( .IN1(n14), .IN2(carry[31]), .Q(SUM[31]) );
  NAND2X0 U24 ( .IN1(A[31]), .IN2(B[31]), .QN(n15) );
  NAND2X0 U25 ( .IN1(A[31]), .IN2(carry[31]), .QN(n16) );
  NAND2X0 U26 ( .IN1(B[31]), .IN2(carry[31]), .QN(n17) );
  NAND3X0 U27 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[32]) );
  XOR3X1 U28 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U29 ( .IN1(A[44]), .IN2(B[44]), .QN(n18) );
  NAND2X0 U30 ( .IN1(A[44]), .IN2(carry[44]), .QN(n19) );
  NAND2X0 U31 ( .IN1(B[44]), .IN2(carry[44]), .QN(n20) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[45]) );
  XOR2X1 U33 ( .IN1(A[45]), .IN2(B[45]), .Q(n21) );
  XOR2X1 U34 ( .IN1(n21), .IN2(carry[45]), .Q(SUM[45]) );
  NAND2X0 U35 ( .IN1(A[45]), .IN2(B[45]), .QN(n22) );
  NAND2X0 U36 ( .IN1(A[45]), .IN2(carry[45]), .QN(n23) );
  NAND2X0 U37 ( .IN1(B[45]), .IN2(carry[45]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[46]) );
  XOR3X1 U39 ( .IN1(carry[43]), .IN2(B[43]), .IN3(A[43]), .Q(SUM[43]) );
  NAND2X0 U40 ( .IN1(A[43]), .IN2(carry[43]), .QN(n25) );
  NAND2X0 U41 ( .IN1(B[43]), .IN2(carry[43]), .QN(n26) );
  NAND2X0 U42 ( .IN1(B[43]), .IN2(A[43]), .QN(n27) );
  NAND3X0 U43 ( .IN1(n25), .IN2(n27), .IN3(n26), .QN(carry[44]) );
  AND2X1 U44 ( .IN1(A[26]), .IN2(B[26]), .Q(n28) );
  XOR2X1 U45 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX2 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  XOR3X1 U1 ( .IN1(carry[38]), .IN2(B[38]), .IN3(A[38]), .Q(SUM[38]) );
  NAND2X1 U2 ( .IN1(A[38]), .IN2(carry[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[38]), .IN2(A[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[39]) );
  XOR3X1 U6 ( .IN1(B[35]), .IN2(A[35]), .IN3(carry[35]), .Q(SUM[35]) );
  NAND2X1 U7 ( .IN1(carry[35]), .IN2(B[35]), .QN(n4) );
  NAND2X1 U8 ( .IN1(A[35]), .IN2(B[35]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[35]), .IN2(carry[35]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[36]) );
  DELLN2X2 U11 ( .INP(carry[48]), .Z(n8) );
  XOR3X1 U12 ( .IN1(B[27]), .IN2(n27), .IN3(A[27]), .Q(SUM[27]) );
  XOR3X1 U13 ( .IN1(A[47]), .IN2(B[47]), .IN3(n7), .Q(SUM[47]) );
  DELLN2X2 U14 ( .INP(carry[47]), .Z(n7) );
  DELLN2X2 U15 ( .INP(carry[45]), .Z(n9) );
  XOR3X2 U16 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  AND2X1 U17 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  NAND2X0 U18 ( .IN1(n27), .IN2(B[27]), .QN(n25) );
  NAND2X0 U19 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U20 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U21 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U22 ( .IN1(n11), .IN2(n12), .IN3(n10), .QN(carry[45]) );
  XOR2X1 U23 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U24 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U25 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U26 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U27 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U28 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U29 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U30 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U31 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U32 ( .IN1(n19), .IN2(n18), .IN3(n17), .QN(carry[48]) );
  XOR2X1 U33 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U34 ( .IN1(n20), .IN2(n8), .Q(SUM[48]) );
  NAND2X0 U35 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U36 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U37 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U38 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[49]) );
  NAND2X0 U39 ( .IN1(A[27]), .IN2(B[27]), .QN(n24) );
  NAND2X0 U40 ( .IN1(n27), .IN2(A[27]), .QN(n26) );
  NAND3X0 U41 ( .IN1(n24), .IN2(n26), .IN3(n25), .QN(carry[28]) );
  XOR2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_4 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N18, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N69, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[4] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n74), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n74), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n13), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n19), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n25), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n31), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n37), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n43), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(combined_b[1]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(n9), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n15), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n21), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n27), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n33), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n39), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n45), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n49), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n65), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n63), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n63), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n63), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n63), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n63), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n63), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n63), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n63), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n63), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n63), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n59), .IN3(N75), .IN4(n57), .IN5(
        product_shift[9]), .IN6(n76), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n59), .IN3(N74), .IN4(n57), .IN5(
        product_shift[8]), .IN6(n56), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n59), .IN3(N73), .IN4(n57), .IN5(
        product_shift[7]), .IN6(n56), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n59), .IN3(N72), .IN4(n57), .IN5(
        product_shift[6]), .IN6(n56), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n59), .IN3(N71), .IN4(n57), .IN5(
        product_shift[5]), .IN6(n56), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n59), .IN3(N116), .IN4(n57), .IN5(
        product_shift[49]), .IN6(n56), .Q(product2[50]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n59), .IN3(N115), .IN4(n57), .IN5(
        product_shift[49]), .IN6(n56), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n59), .IN3(N114), .IN4(n57), .IN5(
        product_shift[48]), .IN6(n56), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n59), .IN3(N113), .IN4(n57), .IN5(
        product_shift[47]), .IN6(n56), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n59), .IN3(N112), .IN4(n57), .IN5(
        product_shift[46]), .IN6(n56), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n59), .IN3(N111), .IN4(n57), .IN5(
        product_shift[45]), .IN6(n56), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n60), .IN3(N110), .IN4(n77), .IN5(
        product_shift[44]), .IN6(n55), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n60), .IN3(N109), .IN4(n77), .IN5(
        product_shift[43]), .IN6(n55), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n60), .IN3(N108), .IN4(n77), .IN5(
        product_shift[42]), .IN6(n55), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n60), .IN3(N107), .IN4(n77), .IN5(
        product_shift[41]), .IN6(n55), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n60), .IN3(N106), .IN4(n77), .IN5(
        product_shift[40]), .IN6(n55), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n60), .IN3(N69), .IN4(n77), .IN5(
        product_shift[3]), .IN6(n55), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n60), .IN3(N105), .IN4(n77), .IN5(
        product_shift[39]), .IN6(n55), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n60), .IN3(N104), .IN4(n77), .IN5(
        product_shift[38]), .IN6(n55), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n60), .IN3(N103), .IN4(n77), .IN5(
        product_shift[37]), .IN6(n55), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n60), .IN3(N102), .IN4(n77), .IN5(
        product_shift[36]), .IN6(n55), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n60), .IN3(N101), .IN4(n77), .IN5(n4), .IN6(
        n55), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n60), .IN3(N100), .IN4(n57), .IN5(n11), .IN6(
        n55), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n61), .IN3(N99), .IN4(n77), .IN5(n17), .IN6(
        n55), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n61), .IN3(N98), .IN4(n58), .IN5(n23), .IN6(
        n76), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n61), .IN3(N97), .IN4(n57), .IN5(n29), .IN6(
        n76), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n61), .IN3(N96), .IN4(n58), .IN5(n35), .IN6(
        n76), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n61), .IN3(N68), .IN4(n58), .IN5(
        product_shift[2]), .IN6(n76), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n61), .IN3(N95), .IN4(n58), .IN5(n41), .IN6(
        n76), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n61), .IN3(N94), .IN4(n58), .IN5(n47), .IN6(
        n76), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n61), .IN3(N93), .IN4(n58), .IN5(n51), .IN6(
        n56), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n61), .IN3(N92), .IN4(n58), .IN5(n53), .IN6(
        n55), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n61), .IN3(N91), .IN4(n58), .IN5(
        product_shift[25]), .IN6(n56), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n61), .IN3(N90), .IN4(n58), .IN5(
        product_shift[24]), .IN6(n55), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n61), .IN3(N89), .IN4(n58), .IN5(
        product_shift[23]), .IN6(n56), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n61), .IN3(N88), .IN4(n77), .IN5(
        product_shift[22]), .IN6(n56), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n62), .IN3(N87), .IN4(n77), .IN5(
        product_shift[21]), .IN6(n76), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n59), .IN3(N86), .IN4(n77), .IN5(
        product_shift[20]), .IN6(n76), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n62), .IN3(N67), .IN4(n58), .IN5(n76), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n62), .IN3(N85), .IN4(n77), .IN5(
        product_shift[19]), .IN6(n76), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n62), .IN3(N84), .IN4(n77), .IN5(
        product_shift[18]), .IN6(n76), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n62), .IN3(N83), .IN4(n77), .IN5(
        product_shift[17]), .IN6(n76), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n62), .IN3(N82), .IN4(n77), .IN5(
        product_shift[16]), .IN6(n76), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n62), .IN3(N81), .IN4(n58), .IN5(
        product_shift[15]), .IN6(n76), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n62), .IN3(N80), .IN4(n57), .IN5(
        product_shift[14]), .IN6(n76), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n62), .IN3(N79), .IN4(n58), .IN5(
        product_shift[13]), .IN6(n76), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n62), .IN3(N78), .IN4(n57), .IN5(
        product_shift[12]), .IN6(n55), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n62), .IN3(N77), .IN4(n58), .IN5(
        product_shift[11]), .IN6(n56), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n62), .IN3(N76), .IN4(n58), .IN5(
        product_shift[10]), .IN6(n56), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n76) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n75), .Q(n77) );
  booth6_4_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:36], n4, 
        n11, n17, n23, n29, n35, n41, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_negative_b[24:9], n9, n15, n21, n27, n33, n39, n45, n49, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, SYNOPSYS_UNCONNECTED__0, N69, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_4_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:36], n4, 
        n11, n17, n23, n29, n35, n41, n47, n51, n53, product_shift[25:0]}), 
        .B({combined_b[24:8], n13, n19, n25, n31, n37, n43, combined_b[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        SYNOPSYS_UNCONNECTED__2, N18, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  INVX0 U3 ( .INP(product_shift[35]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U13 ( .INP(combined_negative_b[8]), .ZN(n5) );
  INVX0 U57 ( .INP(n5), .ZN(n9) );
  INVX0 U60 ( .INP(product_shift[34]), .ZN(n10) );
  INVX0 U61 ( .INP(n10), .ZN(n11) );
  INVX0 U62 ( .INP(combined_b[7]), .ZN(n12) );
  INVX0 U63 ( .INP(n12), .ZN(n13) );
  INVX0 U64 ( .INP(combined_negative_b[7]), .ZN(n14) );
  INVX0 U65 ( .INP(n14), .ZN(n15) );
  INVX0 U66 ( .INP(product_shift[33]), .ZN(n16) );
  INVX0 U67 ( .INP(n16), .ZN(n17) );
  INVX0 U68 ( .INP(combined_b[6]), .ZN(n18) );
  INVX0 U69 ( .INP(n18), .ZN(n19) );
  INVX0 U70 ( .INP(combined_negative_b[6]), .ZN(n20) );
  INVX0 U71 ( .INP(n20), .ZN(n21) );
  INVX0 U72 ( .INP(product_shift[32]), .ZN(n22) );
  INVX0 U73 ( .INP(n22), .ZN(n23) );
  INVX0 U74 ( .INP(combined_b[5]), .ZN(n24) );
  INVX0 U75 ( .INP(n24), .ZN(n25) );
  INVX0 U76 ( .INP(combined_negative_b[5]), .ZN(n26) );
  INVX0 U77 ( .INP(n26), .ZN(n27) );
  INVX0 U78 ( .INP(product_shift[31]), .ZN(n28) );
  INVX0 U79 ( .INP(n28), .ZN(n29) );
  INVX0 U80 ( .INP(combined_b[4]), .ZN(n30) );
  INVX0 U81 ( .INP(n30), .ZN(n31) );
  INVX0 U82 ( .INP(combined_negative_b[4]), .ZN(n32) );
  INVX0 U83 ( .INP(n32), .ZN(n33) );
  INVX0 U84 ( .INP(product_shift[30]), .ZN(n34) );
  INVX0 U85 ( .INP(n34), .ZN(n35) );
  INVX0 U86 ( .INP(combined_b[3]), .ZN(n36) );
  INVX0 U87 ( .INP(n36), .ZN(n37) );
  INVX0 U88 ( .INP(combined_negative_b[3]), .ZN(n38) );
  INVX0 U89 ( .INP(n38), .ZN(n39) );
  INVX0 U90 ( .INP(product_shift[29]), .ZN(n40) );
  INVX0 U91 ( .INP(n40), .ZN(n41) );
  INVX0 U92 ( .INP(combined_b[2]), .ZN(n42) );
  INVX0 U93 ( .INP(n42), .ZN(n43) );
  INVX0 U94 ( .INP(combined_negative_b[2]), .ZN(n44) );
  INVX0 U95 ( .INP(n44), .ZN(n45) );
  INVX0 U96 ( .INP(product_shift[28]), .ZN(n46) );
  INVX0 U97 ( .INP(n46), .ZN(n47) );
  INVX0 U98 ( .INP(combined_negative_b[1]), .ZN(n48) );
  INVX0 U99 ( .INP(n48), .ZN(n49) );
  NBUFFX2 U100 ( .INP(n54), .Z(n63) );
  NBUFFX2 U101 ( .INP(n54), .Z(n64) );
  NBUFFX2 U102 ( .INP(n54), .Z(n65) );
  NBUFFX2 U103 ( .INP(n54), .Z(n66) );
  NBUFFX2 U104 ( .INP(n54), .Z(n67) );
  NBUFFX2 U105 ( .INP(n54), .Z(n68) );
  NBUFFX2 U106 ( .INP(n54), .Z(n69) );
  NBUFFX2 U107 ( .INP(n54), .Z(n71) );
  NBUFFX2 U108 ( .INP(n54), .Z(n72) );
  NBUFFX2 U109 ( .INP(n54), .Z(n73) );
  NBUFFX2 U110 ( .INP(n54), .Z(n74) );
  NBUFFX2 U111 ( .INP(n54), .Z(n70) );
  NBUFFX2 U112 ( .INP(n78), .Z(n61) );
  NBUFFX2 U113 ( .INP(n78), .Z(n60) );
  NBUFFX2 U114 ( .INP(n78), .Z(n59) );
  NBUFFX2 U115 ( .INP(n78), .Z(n62) );
  NBUFFX2 U116 ( .INP(n76), .Z(n55) );
  NBUFFX2 U117 ( .INP(n76), .Z(n56) );
  NBUFFX2 U118 ( .INP(n77), .Z(n57) );
  NBUFFX2 U119 ( .INP(n77), .Z(n58) );
  NBUFFX2 U120 ( .INP(reset), .Z(n54) );
  NOR2X0 U121 ( .IN1(n75), .IN2(product_shift[1]), .QN(n78) );
  INVX0 U122 ( .INP(product_shift[0]), .ZN(n75) );
  INVX0 U124 ( .INP(product_shift[27]), .ZN(n50) );
  INVX0 U125 ( .INP(n50), .ZN(n51) );
  INVX0 U126 ( .INP(product_shift[26]), .ZN(n52) );
  INVX0 U127 ( .INP(n52), .ZN(n53) );
endmodule


module booth6_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n39), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X2 U1 ( .IN1(A[38]), .IN2(B[38]), .IN3(carry[38]), .Q(SUM[38]) );
  NAND2X0 U2 ( .IN1(A[38]), .IN2(B[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(A[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X0 U4 ( .IN1(B[38]), .IN2(carry[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[39]) );
  XOR2X1 U6 ( .IN1(A[39]), .IN2(B[39]), .Q(n4) );
  XOR2X1 U7 ( .IN1(n4), .IN2(carry[39]), .Q(SUM[39]) );
  NAND2X0 U8 ( .IN1(A[39]), .IN2(B[39]), .QN(n5) );
  NAND2X0 U9 ( .IN1(A[39]), .IN2(carry[39]), .QN(n6) );
  NAND2X0 U10 ( .IN1(B[39]), .IN2(carry[39]), .QN(n7) );
  NAND3X0 U11 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[40]) );
  XOR3X2 U12 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  NAND2X0 U13 ( .IN1(A[48]), .IN2(B[48]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[48]), .IN2(carry[48]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[48]), .IN2(carry[48]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[49]) );
  XOR2X1 U17 ( .IN1(A[49]), .IN2(B[49]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X0 U19 ( .IN1(A[49]), .IN2(B[49]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[49]), .IN2(carry[49]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[49]), .IN2(carry[49]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[50]) );
  DELLN2X2 U23 ( .INP(carry[47]), .Z(n15) );
  DELLN2X2 U24 ( .INP(carry[44]), .Z(n16) );
  DELLN2X2 U25 ( .INP(carry[41]), .Z(n17) );
  XOR3X2 U26 ( .IN1(A[46]), .IN2(B[46]), .IN3(carry[46]), .Q(SUM[46]) );
  XOR3X2 U27 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U28 ( .IN1(A[43]), .IN2(B[43]), .IN3(carry[43]), .Q(SUM[43]) );
  NAND2X0 U29 ( .IN1(A[40]), .IN2(B[40]), .QN(n18) );
  NAND2X0 U30 ( .IN1(A[40]), .IN2(carry[40]), .QN(n19) );
  NAND2X0 U31 ( .IN1(B[40]), .IN2(carry[40]), .QN(n20) );
  NAND3X0 U32 ( .IN1(n18), .IN2(n19), .IN3(n20), .QN(carry[41]) );
  XOR2X1 U33 ( .IN1(A[41]), .IN2(B[41]), .Q(n21) );
  XOR2X1 U34 ( .IN1(n21), .IN2(n17), .Q(SUM[41]) );
  NAND2X0 U35 ( .IN1(A[41]), .IN2(B[41]), .QN(n22) );
  NAND2X0 U36 ( .IN1(A[41]), .IN2(carry[41]), .QN(n23) );
  NAND2X0 U37 ( .IN1(B[41]), .IN2(carry[41]), .QN(n24) );
  NAND3X0 U38 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(carry[42]) );
  NAND2X0 U39 ( .IN1(A[43]), .IN2(B[43]), .QN(n25) );
  NAND2X0 U40 ( .IN1(A[43]), .IN2(carry[43]), .QN(n26) );
  NAND2X0 U41 ( .IN1(B[43]), .IN2(carry[43]), .QN(n27) );
  NAND3X0 U42 ( .IN1(n25), .IN2(n26), .IN3(n27), .QN(carry[44]) );
  XOR2X1 U43 ( .IN1(A[44]), .IN2(B[44]), .Q(n28) );
  XOR2X1 U44 ( .IN1(n28), .IN2(n16), .Q(SUM[44]) );
  NAND2X0 U45 ( .IN1(A[44]), .IN2(B[44]), .QN(n29) );
  NAND2X0 U46 ( .IN1(A[44]), .IN2(carry[44]), .QN(n30) );
  NAND2X0 U47 ( .IN1(B[44]), .IN2(carry[44]), .QN(n31) );
  NAND3X0 U48 ( .IN1(n30), .IN2(n31), .IN3(n29), .QN(carry[45]) );
  NAND2X0 U49 ( .IN1(A[46]), .IN2(B[46]), .QN(n32) );
  NAND2X0 U50 ( .IN1(A[46]), .IN2(carry[46]), .QN(n33) );
  NAND2X0 U51 ( .IN1(B[46]), .IN2(carry[46]), .QN(n34) );
  NAND3X0 U52 ( .IN1(n32), .IN2(n33), .IN3(n34), .QN(carry[47]) );
  XOR2X1 U53 ( .IN1(A[47]), .IN2(B[47]), .Q(n35) );
  XOR2X1 U54 ( .IN1(n35), .IN2(n15), .Q(SUM[47]) );
  NAND2X0 U55 ( .IN1(A[47]), .IN2(B[47]), .QN(n36) );
  NAND2X0 U56 ( .IN1(A[47]), .IN2(carry[47]), .QN(n37) );
  NAND2X0 U57 ( .IN1(B[47]), .IN2(carry[47]), .QN(n38) );
  NAND3X0 U58 ( .IN1(n37), .IN2(n38), .IN3(n36), .QN(carry[48]) );
  AND2X1 U59 ( .IN1(A[26]), .IN2(B[26]), .Q(n39) );
  XOR2X1 U60 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(B[34]), .B(n9), .CI(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n24), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  XOR3X1 U1 ( .IN1(carry[42]), .IN2(B[42]), .IN3(A[42]), .Q(SUM[42]) );
  NAND2X0 U2 ( .IN1(A[42]), .IN2(carry[42]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[42]), .IN2(carry[42]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[42]), .IN2(A[42]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[43]) );
  XOR3X1 U6 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U7 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[50]) );
  DELLN2X2 U11 ( .INP(carry[45]), .Z(n7) );
  INVX0 U12 ( .INP(A[34]), .ZN(n8) );
  INVX0 U13 ( .INP(n8), .ZN(n9) );
  XOR3X1 U14 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  XOR3X1 U15 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  NAND2X0 U16 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U17 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U18 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U19 ( .IN1(n10), .IN2(n11), .IN3(n12), .QN(carry[45]) );
  XOR2X1 U20 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U21 ( .IN1(n13), .IN2(n7), .Q(SUM[45]) );
  NAND2X0 U22 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U23 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U24 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U25 ( .IN1(n16), .IN2(n15), .IN3(n14), .QN(carry[46]) );
  NAND2X0 U26 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U27 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U28 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U29 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U30 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U31 ( .IN1(n20), .IN2(carry[48]), .Q(SUM[48]) );
  NAND2X0 U32 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U34 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U35 ( .IN1(n23), .IN2(n22), .IN3(n21), .QN(carry[49]) );
  AND2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(n24) );
  XOR2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_3 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N17, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N68, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product2_o[3] = 1'b0;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n69), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n69), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n69), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n68), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n67), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n66), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[2]  ( .D(product2[2]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[2]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n65), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n65), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n64), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(combined_b[8]), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n15), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n21), .CLK(clk), .RSTB(n64), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n27), .CLK(clk), .RSTB(n63), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n33), .CLK(clk), .RSTB(n63), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n39), .CLK(clk), .RSTB(n63), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n45), .CLK(clk), .RSTB(n63), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n63), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n63), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n62), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n62), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n62), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n4), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n13), .CLK(clk), .RSTB(n62), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n19), .CLK(clk), .RSTB(n61), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n25), .CLK(clk), .RSTB(n61), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n31), .CLK(clk), .RSTB(n61), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n37), .CLK(clk), .RSTB(n61), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n43), .CLK(clk), .RSTB(n61), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n61), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n61), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n60), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n60), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n60), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n60), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n60), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n59), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n58), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n58), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n58), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n58), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n58), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n58), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n58), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n58), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n58), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n58), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n58), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n54), .IN3(N75), .IN4(n72), .IN5(
        product_shift[9]), .IN6(n50), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n54), .IN3(N74), .IN4(n72), .IN5(
        product_shift[8]), .IN6(n71), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n54), .IN3(N73), .IN4(n72), .IN5(
        product_shift[7]), .IN6(n71), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n54), .IN3(N72), .IN4(n72), .IN5(
        product_shift[6]), .IN6(n71), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n54), .IN3(N71), .IN4(n72), .IN5(
        product_shift[5]), .IN6(n71), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(N65), .IN2(n54), .IN3(N116), .IN4(n72), .IN5(
        product_shift[49]), .IN6(n71), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n54), .IN3(N70), .IN4(n72), .IN5(
        product_shift[4]), .IN6(n50), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n54), .IN3(N115), .IN4(n72), .IN5(
        product_shift[49]), .IN6(n51), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n54), .IN3(N114), .IN4(n72), .IN5(
        product_shift[48]), .IN6(n71), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n54), .IN3(N113), .IN4(n72), .IN5(
        product_shift[47]), .IN6(n51), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n54), .IN3(N112), .IN4(n52), .IN5(
        product_shift[46]), .IN6(n71), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n54), .IN3(N111), .IN4(n53), .IN5(
        product_shift[45]), .IN6(n50), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n55), .IN3(N110), .IN4(n72), .IN5(
        product_shift[44]), .IN6(n71), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n55), .IN3(N109), .IN4(n72), .IN5(
        product_shift[43]), .IN6(n71), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n55), .IN3(N108), .IN4(n72), .IN5(
        product_shift[42]), .IN6(n71), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n55), .IN3(N107), .IN4(n72), .IN5(
        product_shift[41]), .IN6(n71), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n55), .IN3(N106), .IN4(n72), .IN5(
        product_shift[40]), .IN6(n71), .Q(product2[40]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n55), .IN3(N105), .IN4(n72), .IN5(
        product_shift[39]), .IN6(n71), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n55), .IN3(N104), .IN4(n72), .IN5(
        product_shift[38]), .IN6(n71), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n55), .IN3(N103), .IN4(n72), .IN5(
        product_shift[37]), .IN6(n71), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n55), .IN3(N102), .IN4(n72), .IN5(
        product_shift[36]), .IN6(n71), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n55), .IN3(N101), .IN4(n72), .IN5(
        product_shift[35]), .IN6(n71), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n55), .IN3(N100), .IN4(n72), .IN5(
        product_shift[34]), .IN6(n71), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n56), .IN3(N99), .IN4(n52), .IN5(n11), .IN6(
        n51), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n56), .IN3(N98), .IN4(n52), .IN5(n17), .IN6(
        n51), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n56), .IN3(N97), .IN4(n52), .IN5(n23), .IN6(
        n51), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n56), .IN3(N96), .IN4(n52), .IN5(n29), .IN6(
        n51), .Q(product2[30]) );
  AO222X1 U35 ( .IN1(N17), .IN2(n56), .IN3(N68), .IN4(n52), .IN5(
        product_shift[2]), .IN6(n51), .Q(product2[2]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n56), .IN3(N95), .IN4(n52), .IN5(n35), .IN6(
        n51), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n56), .IN3(N94), .IN4(n52), .IN5(n41), .IN6(
        n51), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n56), .IN3(N93), .IN4(n52), .IN5(n47), .IN6(
        n51), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n56), .IN3(N92), .IN4(n52), .IN5(n49), .IN6(
        n51), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n56), .IN3(N91), .IN4(n52), .IN5(
        product_shift[25]), .IN6(n51), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n56), .IN3(N90), .IN4(n52), .IN5(
        product_shift[24]), .IN6(n51), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n56), .IN3(N89), .IN4(n52), .IN5(
        product_shift[23]), .IN6(n51), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n57), .IN3(N88), .IN4(n53), .IN5(
        product_shift[22]), .IN6(n51), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n57), .IN3(N87), .IN4(n53), .IN5(
        product_shift[21]), .IN6(n50), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n57), .IN3(N86), .IN4(n53), .IN5(
        product_shift[20]), .IN6(n50), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n57), .IN3(N67), .IN4(n53), .IN5(n50), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n57), .IN3(N85), .IN4(n53), .IN5(
        product_shift[19]), .IN6(n50), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n57), .IN3(N84), .IN4(n53), .IN5(
        product_shift[18]), .IN6(n50), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n57), .IN3(N83), .IN4(n53), .IN5(
        product_shift[17]), .IN6(n50), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n57), .IN3(N82), .IN4(n53), .IN5(
        product_shift[16]), .IN6(n50), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n57), .IN3(N81), .IN4(n53), .IN5(
        product_shift[15]), .IN6(n50), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n57), .IN3(N80), .IN4(n53), .IN5(
        product_shift[14]), .IN6(n50), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n57), .IN3(N79), .IN4(n53), .IN5(
        product_shift[13]), .IN6(n50), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n57), .IN3(N78), .IN4(n53), .IN5(
        product_shift[12]), .IN6(n50), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n55), .IN3(N77), .IN4(n52), .IN5(
        product_shift[11]), .IN6(n50), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n55), .IN3(N76), .IN4(n53), .IN5(
        product_shift[10]), .IN6(n51), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n71) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n70), .Q(n72) );
  booth6_3_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n4, n13, n19, n25, n31, n37, n43, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, SYNOPSYS_UNCONNECTED__0, N68, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_3_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:34], 
        n11, n17, n23, n29, n35, n41, n47, n49, product_shift[25:0]}), .B({
        combined_b[24:8], n9, n15, n21, n27, n33, n39, n45, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        SYNOPSYS_UNCONNECTED__2, N17, N16, SYNOPSYS_UNCONNECTED__3}) );
  NBUFFX2 U3 ( .INP(reset), .Z(n58) );
  NBUFFX2 U4 ( .INP(reset), .Z(n59) );
  NBUFFX2 U24 ( .INP(reset), .Z(n60) );
  NBUFFX2 U57 ( .INP(reset), .Z(n61) );
  NBUFFX2 U60 ( .INP(reset), .Z(n62) );
  NBUFFX2 U61 ( .INP(reset), .Z(n63) );
  NBUFFX2 U62 ( .INP(reset), .Z(n64) );
  NBUFFX2 U63 ( .INP(reset), .Z(n66) );
  NBUFFX2 U64 ( .INP(reset), .Z(n67) );
  NBUFFX2 U65 ( .INP(reset), .Z(n68) );
  NBUFFX2 U66 ( .INP(reset), .Z(n69) );
  INVX0 U67 ( .INP(combined_negative_b[7]), .ZN(n3) );
  INVX0 U68 ( .INP(n3), .ZN(n4) );
  INVX0 U69 ( .INP(combined_b[7]), .ZN(n5) );
  INVX0 U70 ( .INP(n5), .ZN(n9) );
  INVX0 U71 ( .INP(product_shift[33]), .ZN(n10) );
  INVX0 U72 ( .INP(n10), .ZN(n11) );
  INVX0 U73 ( .INP(combined_negative_b[6]), .ZN(n12) );
  INVX0 U74 ( .INP(n12), .ZN(n13) );
  INVX0 U75 ( .INP(combined_b[6]), .ZN(n14) );
  INVX0 U76 ( .INP(n14), .ZN(n15) );
  INVX0 U77 ( .INP(product_shift[32]), .ZN(n16) );
  INVX0 U78 ( .INP(n16), .ZN(n17) );
  INVX0 U79 ( .INP(combined_negative_b[5]), .ZN(n18) );
  INVX0 U80 ( .INP(n18), .ZN(n19) );
  INVX0 U81 ( .INP(combined_b[5]), .ZN(n20) );
  INVX0 U82 ( .INP(n20), .ZN(n21) );
  INVX0 U83 ( .INP(product_shift[31]), .ZN(n22) );
  INVX0 U84 ( .INP(n22), .ZN(n23) );
  INVX0 U85 ( .INP(combined_negative_b[4]), .ZN(n24) );
  INVX0 U86 ( .INP(n24), .ZN(n25) );
  INVX0 U87 ( .INP(combined_b[4]), .ZN(n26) );
  INVX0 U88 ( .INP(n26), .ZN(n27) );
  INVX0 U89 ( .INP(product_shift[30]), .ZN(n28) );
  INVX0 U90 ( .INP(n28), .ZN(n29) );
  INVX0 U91 ( .INP(combined_negative_b[3]), .ZN(n30) );
  INVX0 U92 ( .INP(n30), .ZN(n31) );
  INVX0 U93 ( .INP(combined_b[3]), .ZN(n32) );
  INVX0 U94 ( .INP(n32), .ZN(n33) );
  INVX0 U95 ( .INP(product_shift[29]), .ZN(n34) );
  INVX0 U96 ( .INP(n34), .ZN(n35) );
  INVX0 U97 ( .INP(combined_negative_b[2]), .ZN(n36) );
  INVX0 U98 ( .INP(n36), .ZN(n37) );
  INVX0 U99 ( .INP(combined_b[2]), .ZN(n38) );
  INVX0 U100 ( .INP(n38), .ZN(n39) );
  INVX0 U101 ( .INP(product_shift[28]), .ZN(n40) );
  INVX0 U102 ( .INP(n40), .ZN(n41) );
  INVX0 U103 ( .INP(combined_negative_b[1]), .ZN(n42) );
  INVX0 U104 ( .INP(n42), .ZN(n43) );
  INVX0 U105 ( .INP(combined_b[1]), .ZN(n44) );
  INVX0 U106 ( .INP(n44), .ZN(n45) );
  NBUFFX2 U107 ( .INP(n73), .Z(n57) );
  NBUFFX2 U108 ( .INP(n73), .Z(n56) );
  NBUFFX2 U109 ( .INP(n73), .Z(n54) );
  NBUFFX2 U110 ( .INP(n73), .Z(n55) );
  NBUFFX2 U111 ( .INP(n71), .Z(n50) );
  NBUFFX2 U112 ( .INP(n71), .Z(n51) );
  NBUFFX2 U113 ( .INP(n72), .Z(n53) );
  NBUFFX2 U114 ( .INP(n72), .Z(n52) );
  NBUFFX2 U115 ( .INP(reset), .Z(n65) );
  NOR2X0 U116 ( .IN1(n70), .IN2(product_shift[1]), .QN(n73) );
  INVX0 U117 ( .INP(product_shift[0]), .ZN(n70) );
  INVX0 U119 ( .INP(product_shift[27]), .ZN(n46) );
  INVX0 U120 ( .INP(n46), .ZN(n47) );
  INVX0 U121 ( .INP(product_shift[26]), .ZN(n48) );
  INVX0 U122 ( .INP(n48), .ZN(n49) );
endmodule


module booth6_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[1] = A[1];

  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_34 ( .A(B[34]), .B(A[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n24), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  XOR3X1 U1 ( .IN1(carry[38]), .IN2(B[38]), .IN3(A[38]), .Q(SUM[38]) );
  NAND2X1 U2 ( .IN1(A[38]), .IN2(carry[38]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[38]), .IN2(carry[38]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[38]), .IN2(A[38]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[39]) );
  XOR3X1 U6 ( .IN1(carry[49]), .IN2(B[49]), .IN3(A[49]), .Q(SUM[49]) );
  NAND2X0 U7 ( .IN1(A[49]), .IN2(carry[49]), .QN(n4) );
  NAND2X0 U8 ( .IN1(B[49]), .IN2(carry[49]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[49]), .IN2(A[49]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n6), .IN3(n5), .QN(carry[50]) );
  INVX0 U11 ( .INP(carry[48]), .ZN(n7) );
  INVX0 U12 ( .INP(n7), .ZN(n8) );
  DELLN2X2 U13 ( .INP(carry[45]), .Z(n9) );
  XOR3X2 U14 ( .IN1(A[47]), .IN2(B[47]), .IN3(carry[47]), .Q(SUM[47]) );
  XOR3X2 U15 ( .IN1(A[44]), .IN2(B[44]), .IN3(carry[44]), .Q(SUM[44]) );
  NAND2X0 U16 ( .IN1(A[44]), .IN2(B[44]), .QN(n10) );
  NAND2X0 U17 ( .IN1(A[44]), .IN2(carry[44]), .QN(n11) );
  NAND2X0 U18 ( .IN1(B[44]), .IN2(carry[44]), .QN(n12) );
  NAND3X0 U19 ( .IN1(n12), .IN2(n11), .IN3(n10), .QN(carry[45]) );
  XOR2X1 U20 ( .IN1(A[45]), .IN2(B[45]), .Q(n13) );
  XOR2X1 U21 ( .IN1(n13), .IN2(n9), .Q(SUM[45]) );
  NAND2X0 U22 ( .IN1(A[45]), .IN2(B[45]), .QN(n14) );
  NAND2X0 U23 ( .IN1(A[45]), .IN2(carry[45]), .QN(n15) );
  NAND2X0 U24 ( .IN1(B[45]), .IN2(carry[45]), .QN(n16) );
  NAND3X0 U25 ( .IN1(n14), .IN2(n15), .IN3(n16), .QN(carry[46]) );
  NAND2X0 U26 ( .IN1(A[47]), .IN2(B[47]), .QN(n17) );
  NAND2X0 U27 ( .IN1(A[47]), .IN2(carry[47]), .QN(n18) );
  NAND2X0 U28 ( .IN1(B[47]), .IN2(carry[47]), .QN(n19) );
  NAND3X0 U29 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(carry[48]) );
  XOR2X1 U30 ( .IN1(A[48]), .IN2(B[48]), .Q(n20) );
  XOR2X1 U31 ( .IN1(n20), .IN2(n8), .Q(SUM[48]) );
  NAND2X0 U32 ( .IN1(A[48]), .IN2(B[48]), .QN(n21) );
  NAND2X0 U33 ( .IN1(A[48]), .IN2(carry[48]), .QN(n22) );
  NAND2X0 U34 ( .IN1(B[48]), .IN2(carry[48]), .QN(n23) );
  NAND3X0 U35 ( .IN1(n22), .IN2(n23), .IN3(n21), .QN(carry[49]) );
  AND2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(n24) );
  XOR2X1 U37 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [50:1] carry;
  assign SUM[25] = A[25];
  assign SUM[24] = A[24];
  assign SUM[23] = A[23];
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];
  assign SUM[20] = A[20];
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[1] = A[1];

  FADDX1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FADDX1 U1_35 ( .A(n19), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n28), .CO(carry[28]), .S(SUM[27])
         );
  XOR3X1 U1_50 ( .IN1(A[50]), .IN2(B[50]), .IN3(carry[50]), .Q(SUM[50]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX2 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX2 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX2 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  XOR3X1 U1 ( .IN1(carry[47]), .IN2(B[47]), .IN3(A[47]), .Q(SUM[47]) );
  NAND2X1 U2 ( .IN1(A[47]), .IN2(carry[47]), .QN(n1) );
  NAND2X0 U3 ( .IN1(B[47]), .IN2(carry[47]), .QN(n2) );
  NAND2X1 U4 ( .IN1(B[47]), .IN2(A[47]), .QN(n3) );
  NAND3X0 U5 ( .IN1(n1), .IN2(n3), .IN3(n2), .QN(carry[48]) );
  XOR3X1 U6 ( .IN1(A[45]), .IN2(B[45]), .IN3(carry[45]), .Q(SUM[45]) );
  NAND2X1 U7 ( .IN1(A[45]), .IN2(B[45]), .QN(n4) );
  NAND2X1 U8 ( .IN1(A[45]), .IN2(carry[45]), .QN(n5) );
  NAND2X0 U9 ( .IN1(B[45]), .IN2(carry[45]), .QN(n6) );
  NAND3X0 U10 ( .IN1(n4), .IN2(n5), .IN3(n6), .QN(carry[46]) );
  XOR2X1 U11 ( .IN1(A[46]), .IN2(B[46]), .Q(n7) );
  XOR2X1 U12 ( .IN1(n7), .IN2(carry[46]), .Q(SUM[46]) );
  NAND2X0 U13 ( .IN1(A[46]), .IN2(B[46]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[46]), .IN2(carry[46]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[46]), .IN2(carry[46]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[47]) );
  XOR3X2 U17 ( .IN1(A[39]), .IN2(B[39]), .IN3(carry[39]), .Q(SUM[39]) );
  NAND2X0 U18 ( .IN1(A[39]), .IN2(B[39]), .QN(n11) );
  NAND2X0 U19 ( .IN1(A[39]), .IN2(carry[39]), .QN(n12) );
  NAND2X0 U20 ( .IN1(B[39]), .IN2(carry[39]), .QN(n13) );
  NAND3X0 U21 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(carry[40]) );
  XOR2X1 U22 ( .IN1(A[40]), .IN2(B[40]), .Q(n14) );
  XOR2X1 U23 ( .IN1(n14), .IN2(carry[40]), .Q(SUM[40]) );
  NAND2X0 U24 ( .IN1(A[40]), .IN2(B[40]), .QN(n15) );
  NAND2X0 U25 ( .IN1(A[40]), .IN2(carry[40]), .QN(n16) );
  NAND2X0 U26 ( .IN1(B[40]), .IN2(carry[40]), .QN(n17) );
  NAND3X0 U27 ( .IN1(n15), .IN2(n16), .IN3(n17), .QN(carry[41]) );
  INVX0 U28 ( .INP(A[35]), .ZN(n18) );
  INVX0 U29 ( .INP(n18), .ZN(n19) );
  DELLN2X2 U30 ( .INP(carry[42]), .Z(n20) );
  XOR3X2 U31 ( .IN1(A[41]), .IN2(B[41]), .IN3(carry[41]), .Q(SUM[41]) );
  NAND2X0 U32 ( .IN1(A[41]), .IN2(B[41]), .QN(n21) );
  NAND2X0 U33 ( .IN1(A[41]), .IN2(carry[41]), .QN(n22) );
  NAND2X0 U34 ( .IN1(B[41]), .IN2(carry[41]), .QN(n23) );
  NAND3X0 U35 ( .IN1(n21), .IN2(n22), .IN3(n23), .QN(carry[42]) );
  XOR2X1 U36 ( .IN1(A[42]), .IN2(B[42]), .Q(n24) );
  XOR2X1 U37 ( .IN1(n24), .IN2(n20), .Q(SUM[42]) );
  NAND2X0 U38 ( .IN1(A[42]), .IN2(B[42]), .QN(n25) );
  NAND2X0 U39 ( .IN1(A[42]), .IN2(carry[42]), .QN(n26) );
  NAND2X0 U40 ( .IN1(B[42]), .IN2(carry[42]), .QN(n27) );
  NAND3X0 U41 ( .IN1(n27), .IN2(n26), .IN3(n25), .QN(carry[43]) );
  AND2X1 U42 ( .IN1(A[26]), .IN2(B[26]), .Q(n28) );
  XOR2X1 U43 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_2 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N16, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N67, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, n3, n4, n5, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[1] = product1[2];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n74), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n74), .Q(s2) );
  DFFARX1 \product2_o_reg[50]  ( .D(product2[50]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[50]) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n74), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n73), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[25]) );
  DFFARX1 \product2_o_reg[24]  ( .D(product2[24]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[24]) );
  DFFARX1 \product2_o_reg[23]  ( .D(product2[23]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[23]) );
  DFFARX1 \product2_o_reg[22]  ( .D(product2[22]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[22]) );
  DFFARX1 \product2_o_reg[21]  ( .D(product2[21]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[21]) );
  DFFARX1 \product2_o_reg[20]  ( .D(product2[20]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[20]) );
  DFFARX1 \product2_o_reg[19]  ( .D(product2[19]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[19]) );
  DFFARX1 \product2_o_reg[18]  ( .D(product2[18]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[18]) );
  DFFARX1 \product2_o_reg[17]  ( .D(product2[17]), .CLK(clk), .RSTB(n72), .Q(
        product2_o[17]) );
  DFFARX1 \product2_o_reg[16]  ( .D(product2[16]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[16]) );
  DFFARX1 \product2_o_reg[15]  ( .D(product2[15]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[15]) );
  DFFARX1 \product2_o_reg[14]  ( .D(product2[14]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[14]) );
  DFFARX1 \product2_o_reg[13]  ( .D(product2[13]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[13]) );
  DFFARX1 \product2_o_reg[12]  ( .D(product2[12]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[12]) );
  DFFARX1 \product2_o_reg[11]  ( .D(product2[11]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[11]) );
  DFFARX1 \product2_o_reg[10]  ( .D(product2[10]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[10]) );
  DFFARX1 \product2_o_reg[9]  ( .D(product2[9]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[9]) );
  DFFARX1 \product2_o_reg[8]  ( .D(product2[8]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[8]) );
  DFFARX1 \product2_o_reg[7]  ( .D(product2[7]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[7]) );
  DFFARX1 \product2_o_reg[6]  ( .D(product2[6]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[6]) );
  DFFARX1 \product2_o_reg[5]  ( .D(product2[5]), .CLK(clk), .RSTB(n71), .Q(
        product2_o[5]) );
  DFFARX1 \product2_o_reg[4]  ( .D(product2[4]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[4]) );
  DFFARX1 \product2_o_reg[3]  ( .D(product2[3]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[3]) );
  DFFARX1 \product2_o_reg[1]  ( .D(product2[1]), .CLK(clk), .RSTB(n70), .Q(
        product2_o[1]) );
  DFFARX1 \combined_b2_reg[24]  ( .D(combined_b[24]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[24]) );
  DFFARX1 \combined_b2_reg[23]  ( .D(combined_b[23]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[23]) );
  DFFARX1 \combined_b2_reg[22]  ( .D(combined_b[22]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[22]) );
  DFFARX1 \combined_b2_reg[21]  ( .D(combined_b[21]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[21]) );
  DFFARX1 \combined_b2_reg[20]  ( .D(combined_b[20]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[20]) );
  DFFARX1 \combined_b2_reg[19]  ( .D(combined_b[19]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[19]) );
  DFFARX1 \combined_b2_reg[18]  ( .D(combined_b[18]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[18]) );
  DFFARX1 \combined_b2_reg[17]  ( .D(combined_b[17]), .CLK(clk), .RSTB(n70), 
        .Q(combined_b2[17]) );
  DFFARX1 \combined_b2_reg[16]  ( .D(combined_b[16]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[16]) );
  DFFARX1 \combined_b2_reg[15]  ( .D(combined_b[15]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[15]) );
  DFFARX1 \combined_b2_reg[14]  ( .D(combined_b[14]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[14]) );
  DFFARX1 \combined_b2_reg[13]  ( .D(combined_b[13]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[13]) );
  DFFARX1 \combined_b2_reg[12]  ( .D(combined_b[12]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[12]) );
  DFFARX1 \combined_b2_reg[11]  ( .D(combined_b[11]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[11]) );
  DFFARX1 \combined_b2_reg[10]  ( .D(combined_b[10]), .CLK(clk), .RSTB(n69), 
        .Q(combined_b2[10]) );
  DFFARX1 \combined_b2_reg[9]  ( .D(combined_b[9]), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[9]) );
  DFFARX1 \combined_b2_reg[8]  ( .D(n4), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[8]) );
  DFFARX1 \combined_b2_reg[7]  ( .D(n13), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[7]) );
  DFFARX1 \combined_b2_reg[6]  ( .D(n19), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[6]) );
  DFFARX1 \combined_b2_reg[5]  ( .D(n25), .CLK(clk), .RSTB(n69), .Q(
        combined_b2[5]) );
  DFFARX1 \combined_b2_reg[4]  ( .D(n31), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[4]) );
  DFFARX1 \combined_b2_reg[3]  ( .D(n37), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[3]) );
  DFFARX1 \combined_b2_reg[2]  ( .D(n43), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[2]) );
  DFFARX1 \combined_b2_reg[1]  ( .D(n49), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[1]) );
  DFFARX1 \combined_b2_reg[0]  ( .D(combined_b[0]), .CLK(clk), .RSTB(n68), .Q(
        combined_b2[0]) );
  DFFARX1 \combined_negative_b2_reg[24]  ( .D(combined_negative_b[24]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[24]) );
  DFFARX1 \combined_negative_b2_reg[23]  ( .D(combined_negative_b[23]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[23]) );
  DFFARX1 \combined_negative_b2_reg[22]  ( .D(combined_negative_b[22]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[22]) );
  DFFARX1 \combined_negative_b2_reg[21]  ( .D(combined_negative_b[21]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[21]) );
  DFFARX1 \combined_negative_b2_reg[20]  ( .D(combined_negative_b[20]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[20]) );
  DFFARX1 \combined_negative_b2_reg[19]  ( .D(combined_negative_b[19]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[19]) );
  DFFARX1 \combined_negative_b2_reg[18]  ( .D(combined_negative_b[18]), .CLK(
        clk), .RSTB(n68), .Q(combined_negative_b2[18]) );
  DFFARX1 \combined_negative_b2_reg[17]  ( .D(combined_negative_b[17]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[17]) );
  DFFARX1 \combined_negative_b2_reg[16]  ( .D(combined_negative_b[16]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[16]) );
  DFFARX1 \combined_negative_b2_reg[15]  ( .D(combined_negative_b[15]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[15]) );
  DFFARX1 \combined_negative_b2_reg[14]  ( .D(combined_negative_b[14]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[14]) );
  DFFARX1 \combined_negative_b2_reg[13]  ( .D(combined_negative_b[13]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[13]) );
  DFFARX1 \combined_negative_b2_reg[12]  ( .D(combined_negative_b[12]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[12]) );
  DFFARX1 \combined_negative_b2_reg[11]  ( .D(combined_negative_b[11]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[11]) );
  DFFARX1 \combined_negative_b2_reg[10]  ( .D(combined_negative_b[10]), .CLK(
        clk), .RSTB(n67), .Q(combined_negative_b2[10]) );
  DFFARX1 \combined_negative_b2_reg[9]  ( .D(combined_negative_b[9]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[9]) );
  DFFARX1 \combined_negative_b2_reg[8]  ( .D(combined_negative_b[8]), .CLK(clk), .RSTB(n67), .Q(combined_negative_b2[8]) );
  DFFARX1 \combined_negative_b2_reg[7]  ( .D(n11), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[7]) );
  DFFARX1 \combined_negative_b2_reg[6]  ( .D(n17), .CLK(clk), .RSTB(n67), .Q(
        combined_negative_b2[6]) );
  DFFARX1 \combined_negative_b2_reg[5]  ( .D(n23), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[5]) );
  DFFARX1 \combined_negative_b2_reg[4]  ( .D(n29), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[4]) );
  DFFARX1 \combined_negative_b2_reg[3]  ( .D(n35), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[3]) );
  DFFARX1 \combined_negative_b2_reg[2]  ( .D(n41), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[2]) );
  DFFARX1 \combined_negative_b2_reg[1]  ( .D(n47), .CLK(clk), .RSTB(n66), .Q(
        combined_negative_b2[1]) );
  DFFARX1 \combined_negative_b2_reg[0]  ( .D(combined_negative_b[0]), .CLK(clk), .RSTB(n66), .Q(combined_negative_b2[0]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n66), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n65), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n65), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n65), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n64), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n63), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n63), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n63), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n63), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n63), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n63), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n63), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n63), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n63), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n63), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n63), .Q(add_r2[0])
         );
  AO222X1 U7 ( .IN1(N24), .IN2(n58), .IN3(N75), .IN4(n77), .IN5(
        product_shift[9]), .IN6(n54), .Q(product2[9]) );
  AO222X1 U8 ( .IN1(N23), .IN2(n58), .IN3(N74), .IN4(n77), .IN5(
        product_shift[8]), .IN6(n76), .Q(product2[8]) );
  AO222X1 U9 ( .IN1(N22), .IN2(n58), .IN3(N73), .IN4(n77), .IN5(
        product_shift[7]), .IN6(n76), .Q(product2[7]) );
  AO222X1 U10 ( .IN1(N21), .IN2(n58), .IN3(N72), .IN4(n77), .IN5(
        product_shift[6]), .IN6(n76), .Q(product2[6]) );
  AO222X1 U11 ( .IN1(N20), .IN2(n58), .IN3(N71), .IN4(n77), .IN5(
        product_shift[5]), .IN6(n76), .Q(product2[5]) );
  AO222X1 U12 ( .IN1(n58), .IN2(N65), .IN3(N116), .IN4(n77), .IN5(
        product_shift[49]), .IN6(n76), .Q(product2[50]) );
  AO222X1 U13 ( .IN1(N19), .IN2(n58), .IN3(N70), .IN4(n77), .IN5(
        product_shift[4]), .IN6(n54), .Q(product2[4]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n58), .IN3(N115), .IN4(n77), .IN5(
        product_shift[49]), .IN6(n55), .Q(product2[49]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n58), .IN3(N114), .IN4(n77), .IN5(
        product_shift[48]), .IN6(n76), .Q(product2[48]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n58), .IN3(N113), .IN4(n77), .IN5(
        product_shift[47]), .IN6(n55), .Q(product2[47]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n58), .IN3(N112), .IN4(n56), .IN5(
        product_shift[46]), .IN6(n76), .Q(product2[46]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n58), .IN3(N111), .IN4(n57), .IN5(
        product_shift[45]), .IN6(n76), .Q(product2[45]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n59), .IN3(N110), .IN4(n56), .IN5(
        product_shift[44]), .IN6(n55), .Q(product2[44]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n59), .IN3(N109), .IN4(n56), .IN5(
        product_shift[43]), .IN6(n55), .Q(product2[43]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n59), .IN3(N108), .IN4(n56), .IN5(
        product_shift[42]), .IN6(n55), .Q(product2[42]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n59), .IN3(N107), .IN4(n56), .IN5(
        product_shift[41]), .IN6(n55), .Q(product2[41]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n59), .IN3(N106), .IN4(n56), .IN5(
        product_shift[40]), .IN6(n55), .Q(product2[40]) );
  AO222X1 U24 ( .IN1(N18), .IN2(n59), .IN3(N69), .IN4(n56), .IN5(
        product_shift[3]), .IN6(n55), .Q(product2[3]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n59), .IN3(N105), .IN4(n56), .IN5(
        product_shift[39]), .IN6(n55), .Q(product2[39]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n59), .IN3(N104), .IN4(n56), .IN5(
        product_shift[38]), .IN6(n55), .Q(product2[38]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n59), .IN3(N103), .IN4(n56), .IN5(
        product_shift[37]), .IN6(n55), .Q(product2[37]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n59), .IN3(N102), .IN4(n56), .IN5(
        product_shift[36]), .IN6(n55), .Q(product2[36]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n59), .IN3(N101), .IN4(n56), .IN5(
        product_shift[35]), .IN6(n55), .Q(product2[35]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n59), .IN3(N100), .IN4(n56), .IN5(n9), .IN6(
        n55), .Q(product2[34]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n60), .IN3(N99), .IN4(n77), .IN5(n15), .IN6(
        n55), .Q(product2[33]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n60), .IN3(N98), .IN4(n77), .IN5(n21), .IN6(
        n76), .Q(product2[32]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n60), .IN3(N97), .IN4(n77), .IN5(n27), .IN6(
        n76), .Q(product2[31]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n60), .IN3(N96), .IN4(n77), .IN5(n33), .IN6(
        n76), .Q(product2[30]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n60), .IN3(N95), .IN4(n77), .IN5(n39), .IN6(
        n76), .Q(product2[29]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n60), .IN3(N94), .IN4(n77), .IN5(n45), .IN6(
        n76), .Q(product2[28]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n60), .IN3(N93), .IN4(n77), .IN5(n51), .IN6(
        n76), .Q(product2[27]) );
  AO222X1 U39 ( .IN1(N41), .IN2(n60), .IN3(N92), .IN4(n77), .IN5(n53), .IN6(
        n76), .Q(product2[26]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n60), .IN3(N91), .IN4(n77), .IN5(
        product_shift[25]), .IN6(n76), .Q(product2[25]) );
  AO222X1 U41 ( .IN1(N39), .IN2(n60), .IN3(N90), .IN4(n77), .IN5(
        product_shift[24]), .IN6(n76), .Q(product2[24]) );
  AO222X1 U42 ( .IN1(N38), .IN2(n60), .IN3(N89), .IN4(n77), .IN5(
        product_shift[23]), .IN6(n76), .Q(product2[23]) );
  AO222X1 U43 ( .IN1(N37), .IN2(n61), .IN3(N88), .IN4(n57), .IN5(
        product_shift[22]), .IN6(n54), .Q(product2[22]) );
  AO222X1 U44 ( .IN1(N36), .IN2(n61), .IN3(N87), .IN4(n57), .IN5(
        product_shift[21]), .IN6(n54), .Q(product2[21]) );
  AO222X1 U45 ( .IN1(N35), .IN2(n61), .IN3(N86), .IN4(n57), .IN5(
        product_shift[20]), .IN6(n54), .Q(product2[20]) );
  AO222X1 U46 ( .IN1(N16), .IN2(n61), .IN3(N67), .IN4(n57), .IN5(n54), .IN6(
        product_shift[1]), .Q(product2[1]) );
  AO222X1 U47 ( .IN1(N34), .IN2(n61), .IN3(N85), .IN4(n57), .IN5(
        product_shift[19]), .IN6(n54), .Q(product2[19]) );
  AO222X1 U48 ( .IN1(N33), .IN2(n61), .IN3(N84), .IN4(n57), .IN5(
        product_shift[18]), .IN6(n54), .Q(product2[18]) );
  AO222X1 U49 ( .IN1(N32), .IN2(n61), .IN3(N83), .IN4(n57), .IN5(
        product_shift[17]), .IN6(n54), .Q(product2[17]) );
  AO222X1 U50 ( .IN1(N31), .IN2(n61), .IN3(N82), .IN4(n57), .IN5(
        product_shift[16]), .IN6(n54), .Q(product2[16]) );
  AO222X1 U51 ( .IN1(N30), .IN2(n61), .IN3(N81), .IN4(n57), .IN5(
        product_shift[15]), .IN6(n54), .Q(product2[15]) );
  AO222X1 U52 ( .IN1(N29), .IN2(n61), .IN3(N80), .IN4(n57), .IN5(
        product_shift[14]), .IN6(n54), .Q(product2[14]) );
  AO222X1 U53 ( .IN1(N28), .IN2(n61), .IN3(N79), .IN4(n57), .IN5(
        product_shift[13]), .IN6(n54), .Q(product2[13]) );
  AO222X1 U54 ( .IN1(N27), .IN2(n61), .IN3(N78), .IN4(n57), .IN5(
        product_shift[12]), .IN6(n54), .Q(product2[12]) );
  AO222X1 U55 ( .IN1(N26), .IN2(n62), .IN3(N77), .IN4(n56), .IN5(
        product_shift[11]), .IN6(n54), .Q(product2[11]) );
  AO222X1 U56 ( .IN1(N25), .IN2(n62), .IN3(N76), .IN4(n57), .IN5(
        product_shift[10]), .IN6(n55), .Q(product2[10]) );
  XNOR2X1 U58 ( .IN1(product_shift[0]), .IN2(product_shift[1]), .Q(n76) );
  AND2X1 U59 ( .IN1(product_shift[1]), .IN2(n75), .Q(n77) );
  booth6_2_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:35], n9, 
        n15, n21, n27, n33, n39, n45, n51, n53, product_shift[25:0]}), .B({
        combined_negative_b[24:8], n11, n17, n23, n29, n35, n41, n47, 
        combined_negative_b[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, SYNOPSYS_UNCONNECTED__0, N67, 
        SYNOPSYS_UNCONNECTED__1}) );
  booth6_2_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:35], n9, 
        n15, n21, n27, n33, n39, n45, n51, n53, product_shift[25:0]}), .B({
        combined_b[24:9], n4, n13, n19, n25, n31, n37, n43, n49, combined_b[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        SYNOPSYS_UNCONNECTED__2, N16, SYNOPSYS_UNCONNECTED__3}) );
  NBUFFX2 U3 ( .INP(reset), .Z(n63) );
  NBUFFX2 U4 ( .INP(reset), .Z(n64) );
  NBUFFX2 U35 ( .INP(reset), .Z(n65) );
  NBUFFX2 U57 ( .INP(reset), .Z(n66) );
  NBUFFX2 U60 ( .INP(reset), .Z(n67) );
  NBUFFX2 U61 ( .INP(reset), .Z(n68) );
  NBUFFX2 U62 ( .INP(reset), .Z(n69) );
  NBUFFX2 U63 ( .INP(reset), .Z(n71) );
  NBUFFX2 U64 ( .INP(reset), .Z(n72) );
  NBUFFX2 U65 ( .INP(reset), .Z(n73) );
  NBUFFX2 U66 ( .INP(reset), .Z(n74) );
  INVX0 U67 ( .INP(combined_b[8]), .ZN(n3) );
  INVX0 U68 ( .INP(n3), .ZN(n4) );
  INVX0 U69 ( .INP(product_shift[34]), .ZN(n5) );
  INVX0 U70 ( .INP(n5), .ZN(n9) );
  INVX0 U71 ( .INP(combined_negative_b[7]), .ZN(n10) );
  INVX0 U72 ( .INP(n10), .ZN(n11) );
  INVX0 U73 ( .INP(combined_b[7]), .ZN(n12) );
  INVX0 U74 ( .INP(n12), .ZN(n13) );
  INVX0 U75 ( .INP(product_shift[33]), .ZN(n14) );
  INVX0 U76 ( .INP(n14), .ZN(n15) );
  INVX0 U77 ( .INP(combined_negative_b[6]), .ZN(n16) );
  INVX0 U78 ( .INP(n16), .ZN(n17) );
  INVX0 U79 ( .INP(combined_b[6]), .ZN(n18) );
  INVX0 U80 ( .INP(n18), .ZN(n19) );
  INVX0 U81 ( .INP(product_shift[32]), .ZN(n20) );
  INVX0 U82 ( .INP(n20), .ZN(n21) );
  INVX0 U83 ( .INP(combined_negative_b[5]), .ZN(n22) );
  INVX0 U84 ( .INP(n22), .ZN(n23) );
  INVX0 U85 ( .INP(combined_b[5]), .ZN(n24) );
  INVX0 U86 ( .INP(n24), .ZN(n25) );
  INVX0 U87 ( .INP(product_shift[31]), .ZN(n26) );
  INVX0 U88 ( .INP(n26), .ZN(n27) );
  INVX0 U89 ( .INP(combined_negative_b[4]), .ZN(n28) );
  INVX0 U90 ( .INP(n28), .ZN(n29) );
  INVX0 U91 ( .INP(combined_b[4]), .ZN(n30) );
  INVX0 U92 ( .INP(n30), .ZN(n31) );
  INVX0 U93 ( .INP(product_shift[30]), .ZN(n32) );
  INVX0 U94 ( .INP(n32), .ZN(n33) );
  INVX0 U95 ( .INP(combined_negative_b[3]), .ZN(n34) );
  INVX0 U96 ( .INP(n34), .ZN(n35) );
  INVX0 U97 ( .INP(combined_b[3]), .ZN(n36) );
  INVX0 U98 ( .INP(n36), .ZN(n37) );
  INVX0 U99 ( .INP(product_shift[29]), .ZN(n38) );
  INVX0 U100 ( .INP(n38), .ZN(n39) );
  INVX0 U101 ( .INP(combined_negative_b[2]), .ZN(n40) );
  INVX0 U102 ( .INP(n40), .ZN(n41) );
  INVX0 U103 ( .INP(combined_b[2]), .ZN(n42) );
  INVX0 U104 ( .INP(n42), .ZN(n43) );
  INVX0 U105 ( .INP(product_shift[28]), .ZN(n44) );
  INVX0 U106 ( .INP(n44), .ZN(n45) );
  INVX0 U107 ( .INP(combined_negative_b[1]), .ZN(n46) );
  INVX0 U108 ( .INP(n46), .ZN(n47) );
  INVX0 U109 ( .INP(combined_b[1]), .ZN(n48) );
  INVX0 U110 ( .INP(n48), .ZN(n49) );
  NBUFFX2 U111 ( .INP(n78), .Z(n61) );
  NBUFFX2 U112 ( .INP(n78), .Z(n59) );
  NBUFFX2 U113 ( .INP(n78), .Z(n58) );
  NBUFFX2 U114 ( .INP(n78), .Z(n60) );
  NBUFFX2 U115 ( .INP(n78), .Z(n62) );
  NBUFFX2 U116 ( .INP(n76), .Z(n54) );
  NBUFFX2 U117 ( .INP(n76), .Z(n55) );
  NBUFFX2 U118 ( .INP(n77), .Z(n57) );
  NBUFFX2 U119 ( .INP(n77), .Z(n56) );
  NBUFFX2 U120 ( .INP(reset), .Z(n70) );
  NOR2X0 U121 ( .IN1(n75), .IN2(product_shift[1]), .QN(n78) );
  INVX0 U122 ( .INP(product_shift[0]), .ZN(n75) );
  INVX0 U123 ( .INP(product_shift[27]), .ZN(n50) );
  INVX0 U124 ( .INP(n50), .ZN(n51) );
  INVX0 U125 ( .INP(product_shift[26]), .ZN(n52) );
  INVX0 U126 ( .INP(n52), .ZN(n53) );
endmodule


module booth6_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [50:1] carry;
  assign SUM[25] = A[25];

  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FADDX1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n1), .CO(carry[28]), .S(SUM[27]) );
  XOR3X1 U1_49 ( .IN1(A[49]), .IN2(B[49]), .IN3(carry[49]), .Q(SUM[49]) );
  AND2X1 U1 ( .IN1(A[26]), .IN2(B[26]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [50:0] A;
  input [50:0] B;
  output [50:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [50:1] carry;
  assign SUM[25] = A[25];

  FADDX1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(n16), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_31 ( .A(A[31]), .B(n18), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(n20), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(n22), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(n24), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(n26), .CI(n27), .CO(carry[28]), .S(SUM[27]) );
  XOR3X1 U1_49 ( .IN1(A[49]), .IN2(B[49]), .IN3(carry[49]), .Q(SUM[49]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FADDX1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FADDX1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FADDX1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  XOR3X1 U1 ( .IN1(A[34]), .IN2(B[34]), .IN3(carry[34]), .Q(SUM[34]) );
  XOR3X1 U2 ( .IN1(A[41]), .IN2(B[41]), .IN3(carry[41]), .Q(SUM[41]) );
  NAND2X0 U3 ( .IN1(A[41]), .IN2(B[41]), .QN(n1) );
  NAND2X0 U4 ( .IN1(A[41]), .IN2(carry[41]), .QN(n2) );
  NAND2X0 U5 ( .IN1(B[41]), .IN2(carry[41]), .QN(n3) );
  NAND3X0 U6 ( .IN1(n1), .IN2(n2), .IN3(n3), .QN(carry[42]) );
  XOR2X1 U7 ( .IN1(A[42]), .IN2(B[42]), .Q(n4) );
  XOR2X1 U8 ( .IN1(n4), .IN2(carry[42]), .Q(SUM[42]) );
  NAND2X0 U9 ( .IN1(A[42]), .IN2(B[42]), .QN(n5) );
  NAND2X0 U10 ( .IN1(A[42]), .IN2(carry[42]), .QN(n6) );
  NAND2X0 U11 ( .IN1(B[42]), .IN2(carry[42]), .QN(n7) );
  NAND3X0 U12 ( .IN1(n5), .IN2(n6), .IN3(n7), .QN(carry[43]) );
  NAND2X0 U13 ( .IN1(A[34]), .IN2(B[34]), .QN(n8) );
  NAND2X0 U14 ( .IN1(A[34]), .IN2(carry[34]), .QN(n9) );
  NAND2X0 U15 ( .IN1(B[34]), .IN2(carry[34]), .QN(n10) );
  NAND3X0 U16 ( .IN1(n8), .IN2(n9), .IN3(n10), .QN(carry[35]) );
  XOR2X1 U17 ( .IN1(A[35]), .IN2(B[35]), .Q(n11) );
  XOR2X1 U18 ( .IN1(n11), .IN2(carry[35]), .Q(SUM[35]) );
  NAND2X0 U19 ( .IN1(A[35]), .IN2(B[35]), .QN(n12) );
  NAND2X0 U20 ( .IN1(A[35]), .IN2(carry[35]), .QN(n13) );
  NAND2X0 U21 ( .IN1(B[35]), .IN2(carry[35]), .QN(n14) );
  NAND3X0 U22 ( .IN1(n12), .IN2(n13), .IN3(n14), .QN(carry[36]) );
  INVX0 U23 ( .INP(B[32]), .ZN(n15) );
  INVX0 U24 ( .INP(n15), .ZN(n16) );
  INVX0 U25 ( .INP(B[31]), .ZN(n17) );
  INVX0 U26 ( .INP(n17), .ZN(n18) );
  INVX0 U27 ( .INP(B[30]), .ZN(n19) );
  INVX0 U28 ( .INP(n19), .ZN(n20) );
  INVX0 U29 ( .INP(B[29]), .ZN(n21) );
  INVX0 U30 ( .INP(n21), .ZN(n22) );
  INVX0 U31 ( .INP(B[28]), .ZN(n23) );
  INVX0 U32 ( .INP(n23), .ZN(n24) );
  INVX0 U33 ( .INP(B[27]), .ZN(n25) );
  INVX0 U34 ( .INP(n25), .ZN(n26) );
  AND2X1 U35 ( .IN1(A[26]), .IN2(B[26]), .Q(n27) );
  XOR2X1 U36 ( .IN1(A[26]), .IN2(B[26]), .Q(SUM[26]) );
endmodule


module booth6_1 ( clk, reset, product1, combined_b, combined_negative_b, 
        product2_o, combined_b2, combined_negative_b2, new_exponent, 
        new_exponent2, new_sign, new_sign2, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [50:0] product1;
  input [24:0] combined_b;
  input [24:0] combined_negative_b;
  output [50:0] product2_o;
  output [24:0] combined_b2;
  output [24:0] combined_negative_b2;
  input [8:0] new_exponent;
  output [8:0] new_exponent2;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output new_sign2, add_exception_2, s2;
  wire   N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, n4, n5,
         n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39;
  wire   [50:0] product2;
  wire   [50:0] product_shift;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51;
  assign product_shift[49] = product1[50];
  assign product_shift[48] = product1[49];
  assign product_shift[47] = product1[48];
  assign product_shift[46] = product1[47];
  assign product_shift[45] = product1[46];
  assign product_shift[44] = product1[45];
  assign product_shift[43] = product1[44];
  assign product_shift[42] = product1[43];
  assign product_shift[41] = product1[42];
  assign product_shift[40] = product1[41];
  assign product_shift[39] = product1[40];
  assign product_shift[38] = product1[39];
  assign product_shift[37] = product1[38];
  assign product_shift[36] = product1[37];
  assign product_shift[35] = product1[36];
  assign product_shift[34] = product1[35];
  assign product_shift[33] = product1[34];
  assign product_shift[32] = product1[33];
  assign product_shift[31] = product1[32];
  assign product_shift[30] = product1[31];
  assign product_shift[29] = product1[30];
  assign product_shift[28] = product1[29];
  assign product_shift[27] = product1[28];
  assign product_shift[26] = product1[27];
  assign product_shift[25] = product1[26];
  assign product_shift[24] = product1[25];
  assign product_shift[23] = product1[24];
  assign product_shift[22] = product1[23];
  assign product_shift[21] = product1[22];
  assign product_shift[20] = product1[21];
  assign product_shift[19] = product1[20];
  assign product_shift[18] = product1[19];
  assign product_shift[17] = product1[18];
  assign product_shift[16] = product1[17];
  assign product_shift[15] = product1[16];
  assign product_shift[14] = product1[15];
  assign product_shift[13] = product1[14];
  assign product_shift[12] = product1[13];
  assign product_shift[11] = product1[12];
  assign product_shift[10] = product1[11];
  assign product_shift[9] = product1[10];
  assign product_shift[8] = product1[9];
  assign product_shift[7] = product1[8];
  assign product_shift[6] = product1[7];
  assign product_shift[5] = product1[6];
  assign product_shift[4] = product1[5];
  assign product_shift[3] = product1[4];
  assign product_shift[2] = product1[3];
  assign product_shift[0] = product1[1];

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n36), 
        .Q(add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n36), .Q(s2) );
  DFFARX1 \product2_o_reg[49]  ( .D(product2[49]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[49]) );
  DFFARX1 \product2_o_reg[48]  ( .D(product2[48]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[48]) );
  DFFARX1 \product2_o_reg[47]  ( .D(product2[47]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[47]) );
  DFFARX1 \product2_o_reg[46]  ( .D(product2[46]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[46]) );
  DFFARX1 \product2_o_reg[45]  ( .D(product2[45]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[45]) );
  DFFARX1 \product2_o_reg[44]  ( .D(product2[44]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[44]) );
  DFFARX1 \product2_o_reg[43]  ( .D(product2[43]), .CLK(clk), .RSTB(n36), .Q(
        product2_o[43]) );
  DFFARX1 \product2_o_reg[42]  ( .D(product2[42]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[42]) );
  DFFARX1 \product2_o_reg[41]  ( .D(product2[41]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[41]) );
  DFFARX1 \product2_o_reg[40]  ( .D(product2[40]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[40]) );
  DFFARX1 \product2_o_reg[39]  ( .D(product2[39]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[39]) );
  DFFARX1 \product2_o_reg[38]  ( .D(product2[38]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[38]) );
  DFFARX1 \product2_o_reg[37]  ( .D(product2[37]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[37]) );
  DFFARX1 \product2_o_reg[36]  ( .D(product2[36]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[36]) );
  DFFARX1 \product2_o_reg[35]  ( .D(product2[35]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[35]) );
  DFFARX1 \product2_o_reg[34]  ( .D(product2[34]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[34]) );
  DFFARX1 \product2_o_reg[33]  ( .D(product2[33]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[33]) );
  DFFARX1 \product2_o_reg[32]  ( .D(product2[32]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[32]) );
  DFFARX1 \product2_o_reg[31]  ( .D(product2[31]), .CLK(clk), .RSTB(n35), .Q(
        product2_o[31]) );
  DFFARX1 \product2_o_reg[30]  ( .D(product2[30]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[30]) );
  DFFARX1 \product2_o_reg[29]  ( .D(product2[29]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[29]) );
  DFFARX1 \product2_o_reg[28]  ( .D(product2[28]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[28]) );
  DFFARX1 \product2_o_reg[27]  ( .D(product2[27]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[27]) );
  DFFARX1 \product2_o_reg[26]  ( .D(product2[26]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[26]) );
  DFFARX1 \product2_o_reg[25]  ( .D(product2[25]), .CLK(clk), .RSTB(n34), .Q(
        product2_o[25]) );
  DFFARX1 \new_exponent2_reg[8]  ( .D(new_exponent[8]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[8]) );
  DFFARX1 \new_exponent2_reg[7]  ( .D(new_exponent[7]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[7]) );
  DFFARX1 \new_exponent2_reg[6]  ( .D(new_exponent[6]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[6]) );
  DFFARX1 \new_exponent2_reg[5]  ( .D(new_exponent[5]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[5]) );
  DFFARX1 \new_exponent2_reg[4]  ( .D(new_exponent[4]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[4]) );
  DFFARX1 \new_exponent2_reg[3]  ( .D(new_exponent[3]), .CLK(clk), .RSTB(n34), 
        .Q(new_exponent2[3]) );
  DFFARX1 \new_exponent2_reg[2]  ( .D(new_exponent[2]), .CLK(clk), .RSTB(n33), 
        .Q(new_exponent2[2]) );
  DFFARX1 \new_exponent2_reg[1]  ( .D(new_exponent[1]), .CLK(clk), .RSTB(n33), 
        .Q(new_exponent2[1]) );
  DFFARX1 \new_exponent2_reg[0]  ( .D(new_exponent[0]), .CLK(clk), .RSTB(n33), 
        .Q(new_exponent2[0]) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n33), .Q(new_sign2)
         );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n33), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n32), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n31), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n31), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n31), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n31), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n31), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n31), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n31), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n31), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n31), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n31), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n31), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n31), .Q(add_r2[0])
         );
  booth6_1_DW01_add_0 add_89 ( .A({product_shift[49], product_shift[49:35], n5, 
        n9, n11, n13, n15, n17, n19, n21, n23, product_shift[25:2], 1'b0, 
        product_shift[0]}), .B({combined_negative_b, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25}) );
  booth6_1_DW01_add_1 add_82 ( .A({product_shift[49], product_shift[49:35], n5, 
        n9, n11, n13, n15, n17, n19, n21, n23, product_shift[25:2], 1'b0, 
        product_shift[0]}), .B({combined_b, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__26, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51}) );
  AO222X1 U39 ( .IN1(N41), .IN2(n30), .IN3(N92), .IN4(1'b0), .IN5(n23), .IN6(
        n25), .Q(product2[26]) );
  AO222X1 U38 ( .IN1(N42), .IN2(n30), .IN3(N93), .IN4(1'b0), .IN5(n21), .IN6(
        n25), .Q(product2[27]) );
  AO222X1 U37 ( .IN1(N43), .IN2(n30), .IN3(N94), .IN4(1'b0), .IN5(n19), .IN6(
        n25), .Q(product2[28]) );
  AO222X1 U36 ( .IN1(N44), .IN2(n30), .IN3(N95), .IN4(1'b0), .IN5(n17), .IN6(
        n25), .Q(product2[29]) );
  AO222X1 U34 ( .IN1(N45), .IN2(n30), .IN3(N96), .IN4(1'b0), .IN5(n15), .IN6(
        n25), .Q(product2[30]) );
  AO222X1 U33 ( .IN1(N46), .IN2(n30), .IN3(N97), .IN4(1'b0), .IN5(n13), .IN6(
        n25), .Q(product2[31]) );
  AO222X1 U32 ( .IN1(N47), .IN2(n30), .IN3(N98), .IN4(1'b0), .IN5(n11), .IN6(
        n25), .Q(product2[32]) );
  AO222X1 U31 ( .IN1(N48), .IN2(n30), .IN3(N99), .IN4(1'b0), .IN5(n9), .IN6(
        n25), .Q(product2[33]) );
  AO222X1 U30 ( .IN1(N49), .IN2(n30), .IN3(N100), .IN4(1'b0), .IN5(n5), .IN6(
        n25), .Q(product2[34]) );
  AO222X1 U29 ( .IN1(N50), .IN2(n30), .IN3(N101), .IN4(1'b0), .IN5(
        product_shift[35]), .IN6(n25), .Q(product2[35]) );
  AO222X1 U28 ( .IN1(N51), .IN2(n30), .IN3(N102), .IN4(1'b0), .IN5(
        product_shift[36]), .IN6(n25), .Q(product2[36]) );
  AO222X1 U27 ( .IN1(N52), .IN2(n30), .IN3(N103), .IN4(1'b0), .IN5(
        product_shift[37]), .IN6(n25), .Q(product2[37]) );
  AO222X1 U40 ( .IN1(N40), .IN2(n30), .IN3(N91), .IN4(1'b0), .IN5(
        product_shift[25]), .IN6(n25), .Q(product2[25]) );
  AO222X1 U26 ( .IN1(N53), .IN2(n29), .IN3(N104), .IN4(1'b0), .IN5(
        product_shift[38]), .IN6(n24), .Q(product2[38]) );
  AO222X1 U25 ( .IN1(N54), .IN2(n29), .IN3(N105), .IN4(1'b0), .IN5(
        product_shift[39]), .IN6(n24), .Q(product2[39]) );
  AO222X1 U23 ( .IN1(N55), .IN2(n29), .IN3(N106), .IN4(1'b0), .IN5(
        product_shift[40]), .IN6(n24), .Q(product2[40]) );
  AO222X1 U22 ( .IN1(N56), .IN2(n29), .IN3(N107), .IN4(1'b0), .IN5(
        product_shift[41]), .IN6(n24), .Q(product2[41]) );
  AO222X1 U21 ( .IN1(N57), .IN2(n29), .IN3(N108), .IN4(1'b0), .IN5(
        product_shift[42]), .IN6(n24), .Q(product2[42]) );
  AO222X1 U20 ( .IN1(N58), .IN2(n29), .IN3(N109), .IN4(1'b0), .IN5(
        product_shift[43]), .IN6(n24), .Q(product2[43]) );
  AO222X1 U19 ( .IN1(N59), .IN2(n29), .IN3(N110), .IN4(1'b0), .IN5(
        product_shift[44]), .IN6(n24), .Q(product2[44]) );
  AO222X1 U18 ( .IN1(N60), .IN2(n29), .IN3(N111), .IN4(1'b0), .IN5(
        product_shift[45]), .IN6(n24), .Q(product2[45]) );
  AO222X1 U17 ( .IN1(N61), .IN2(n29), .IN3(N112), .IN4(1'b0), .IN5(
        product_shift[46]), .IN6(n24), .Q(product2[46]) );
  AO222X1 U16 ( .IN1(N62), .IN2(n29), .IN3(N113), .IN4(1'b0), .IN5(
        product_shift[47]), .IN6(n24), .Q(product2[47]) );
  AO222X1 U15 ( .IN1(N63), .IN2(n29), .IN3(N114), .IN4(1'b0), .IN5(
        product_shift[48]), .IN6(n24), .Q(product2[48]) );
  AO222X1 U14 ( .IN1(N64), .IN2(n29), .IN3(N115), .IN4(1'b0), .IN5(
        product_shift[49]), .IN6(n24), .Q(product2[49]) );
  INVX1 U3 ( .INP(product_shift[0]), .ZN(n38) );
  NOR2X0 U4 ( .IN1(n37), .IN2(1'b0), .QN(n39) );
  INVX0 U8 ( .INP(product_shift[34]), .ZN(n4) );
  INVX0 U9 ( .INP(n4), .ZN(n5) );
  INVX0 U10 ( .INP(product_shift[33]), .ZN(n7) );
  INVX0 U11 ( .INP(n7), .ZN(n9) );
  INVX0 U12 ( .INP(product_shift[32]), .ZN(n10) );
  INVX0 U13 ( .INP(n10), .ZN(n11) );
  INVX0 U24 ( .INP(product_shift[31]), .ZN(n12) );
  INVX0 U35 ( .INP(n12), .ZN(n13) );
  INVX0 U41 ( .INP(product_shift[30]), .ZN(n14) );
  INVX0 U42 ( .INP(n14), .ZN(n15) );
  INVX0 U43 ( .INP(product_shift[29]), .ZN(n16) );
  INVX0 U44 ( .INP(n16), .ZN(n17) );
  INVX0 U45 ( .INP(product_shift[28]), .ZN(n18) );
  INVX0 U46 ( .INP(n18), .ZN(n19) );
  INVX0 U47 ( .INP(product_shift[27]), .ZN(n20) );
  INVX0 U48 ( .INP(n20), .ZN(n21) );
  NBUFFX2 U49 ( .INP(n38), .Z(n25) );
  NBUFFX2 U50 ( .INP(n38), .Z(n24) );
  NBUFFX2 U51 ( .INP(n39), .Z(n30) );
  NBUFFX2 U52 ( .INP(n39), .Z(n29) );
  NBUFFX2 U53 ( .INP(reset), .Z(n31) );
  NBUFFX2 U54 ( .INP(reset), .Z(n32) );
  NBUFFX2 U55 ( .INP(reset), .Z(n33) );
  NBUFFX2 U56 ( .INP(reset), .Z(n34) );
  NBUFFX2 U57 ( .INP(reset), .Z(n35) );
  NBUFFX2 U58 ( .INP(reset), .Z(n36) );
  INVX0 U59 ( .INP(product_shift[0]), .ZN(n37) );
  INVX0 U63 ( .INP(product_shift[26]), .ZN(n22) );
  INVX0 U64 ( .INP(n22), .ZN(n23) );
endmodule


module normalize1_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(SUM[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module normalize1_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[8]), .IN2(A[8]), .Q(SUM[8]) );
endmodule


module normalize1 ( clk, reset, product, new_exponent, updated_exponent_o, 
        updated_product_o, exception_o, new_sign, new_sign2, add_r, 
        add_exception_1, add_r2, add_exception_2, s, s2 );
  input [50:0] product;
  input [8:0] new_exponent;
  output [8:0] updated_exponent_o;
  output [24:0] updated_product_o;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, add_exception_1, s;
  output exception_o, new_sign2, add_exception_2, s2;
  wire   N7, N13, N14, N15, N16, N17, N18, N19, N20, N21, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31;
  wire   [8:0] updated_exponent;
  wire   [24:0] updated_product;

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n8), .Q(
        add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n8), .Q(s2) );
  DFFARX1 \updated_exponent_o_reg[8]  ( .D(updated_exponent[8]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[8]) );
  DFFARX1 \updated_exponent_o_reg[7]  ( .D(updated_exponent[7]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[7]) );
  DFFARX1 \updated_exponent_o_reg[6]  ( .D(updated_exponent[6]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[6]) );
  DFFARX1 \updated_exponent_o_reg[5]  ( .D(updated_exponent[5]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[5]) );
  DFFARX1 \updated_exponent_o_reg[4]  ( .D(updated_exponent[4]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[4]) );
  DFFARX1 \updated_exponent_o_reg[3]  ( .D(updated_exponent[3]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[3]) );
  DFFARX1 \updated_exponent_o_reg[2]  ( .D(updated_exponent[2]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[2]) );
  DFFARX1 \updated_exponent_o_reg[1]  ( .D(updated_exponent[1]), .CLK(clk), 
        .RSTB(n8), .Q(updated_exponent_o[1]) );
  DFFARX1 \updated_exponent_o_reg[0]  ( .D(updated_exponent[0]), .CLK(clk), 
        .RSTB(n7), .Q(updated_exponent_o[0]) );
  DFFARX1 \updated_product_o_reg[24]  ( .D(updated_product[24]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[24]) );
  DFFARX1 \updated_product_o_reg[23]  ( .D(updated_product[23]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[23]) );
  DFFARX1 \updated_product_o_reg[22]  ( .D(updated_product[22]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[22]) );
  DFFARX1 \updated_product_o_reg[21]  ( .D(updated_product[21]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[21]) );
  DFFARX1 \updated_product_o_reg[20]  ( .D(updated_product[20]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[20]) );
  DFFARX1 \updated_product_o_reg[19]  ( .D(updated_product[19]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[19]) );
  DFFARX1 \updated_product_o_reg[18]  ( .D(updated_product[18]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[18]) );
  DFFARX1 \updated_product_o_reg[17]  ( .D(updated_product[17]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[17]) );
  DFFARX1 \updated_product_o_reg[16]  ( .D(updated_product[16]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[16]) );
  DFFARX1 \updated_product_o_reg[15]  ( .D(updated_product[15]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[15]) );
  DFFARX1 \updated_product_o_reg[14]  ( .D(updated_product[14]), .CLK(clk), 
        .RSTB(n7), .Q(updated_product_o[14]) );
  DFFARX1 \updated_product_o_reg[13]  ( .D(updated_product[13]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[13]) );
  DFFARX1 \updated_product_o_reg[12]  ( .D(updated_product[12]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[12]) );
  DFFARX1 \updated_product_o_reg[11]  ( .D(updated_product[11]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[11]) );
  DFFARX1 \updated_product_o_reg[10]  ( .D(updated_product[10]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[10]) );
  DFFARX1 \updated_product_o_reg[9]  ( .D(updated_product[9]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[9]) );
  DFFARX1 \updated_product_o_reg[8]  ( .D(updated_product[8]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[8]) );
  DFFARX1 \updated_product_o_reg[7]  ( .D(updated_product[7]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[7]) );
  DFFARX1 \updated_product_o_reg[6]  ( .D(updated_product[6]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[6]) );
  DFFARX1 \updated_product_o_reg[5]  ( .D(updated_product[5]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[5]) );
  DFFARX1 \updated_product_o_reg[4]  ( .D(updated_product[4]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[4]) );
  DFFARX1 \updated_product_o_reg[3]  ( .D(updated_product[3]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[3]) );
  DFFARX1 \updated_product_o_reg[2]  ( .D(updated_product[2]), .CLK(clk), 
        .RSTB(n6), .Q(updated_product_o[2]) );
  DFFARX1 \updated_product_o_reg[1]  ( .D(updated_product[1]), .CLK(clk), 
        .RSTB(n5), .Q(updated_product_o[1]) );
  DFFARX1 \updated_product_o_reg[0]  ( .D(updated_product[0]), .CLK(clk), 
        .RSTB(n5), .Q(updated_product_o[0]) );
  DFFARX1 exception_o_reg ( .D(N7), .CLK(clk), .RSTB(n5), .Q(exception_o) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n5), .Q(new_sign2) );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n3), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n3), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n3), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n3), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n3), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n3), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n3), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n3), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n3), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n3), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n3), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n3), .Q(add_r2[0])
         );
  normalize1_DW01_inc_0 add_95 ( .A({1'b0, product[49:26]}), .SUM({N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23}) );
  normalize1_DW01_inc_1 r66 ( .A(new_exponent), .SUM({N21, N20, N19, N18, N17, 
        N16, N15, N14, N13}) );
  NOR2X0 U3 ( .IN1(n14), .IN2(N7), .QN(n2) );
  OR2X1 U4 ( .IN1(n9), .IN2(n10), .Q(n12) );
  NBUFFX2 U5 ( .INP(reset), .Z(n3) );
  NBUFFX2 U6 ( .INP(reset), .Z(n4) );
  NBUFFX2 U8 ( .INP(reset), .Z(n5) );
  NBUFFX2 U9 ( .INP(reset), .Z(n6) );
  NBUFFX2 U10 ( .INP(reset), .Z(n7) );
  NBUFFX2 U11 ( .INP(reset), .Z(n8) );
  AO222X1 U12 ( .IN1(N32), .IN2(n9), .IN3(product[35]), .IN4(n10), .IN5(
        product[34]), .IN6(n11), .Q(updated_product[9]) );
  AO222X1 U13 ( .IN1(N31), .IN2(n9), .IN3(product[34]), .IN4(n10), .IN5(
        product[33]), .IN6(n2), .Q(updated_product[8]) );
  AO222X1 U14 ( .IN1(N30), .IN2(n9), .IN3(product[33]), .IN4(n10), .IN5(
        product[32]), .IN6(n2), .Q(updated_product[7]) );
  AO222X1 U15 ( .IN1(N29), .IN2(n9), .IN3(product[32]), .IN4(n10), .IN5(
        product[31]), .IN6(n2), .Q(updated_product[6]) );
  AO222X1 U16 ( .IN1(N28), .IN2(n9), .IN3(product[31]), .IN4(n10), .IN5(
        product[30]), .IN6(n2), .Q(updated_product[5]) );
  AO222X1 U17 ( .IN1(N27), .IN2(n9), .IN3(product[30]), .IN4(n10), .IN5(
        product[29]), .IN6(n2), .Q(updated_product[4]) );
  AO222X1 U18 ( .IN1(N26), .IN2(n9), .IN3(product[29]), .IN4(n10), .IN5(
        product[28]), .IN6(n2), .Q(updated_product[3]) );
  AO222X1 U19 ( .IN1(N25), .IN2(n9), .IN3(product[28]), .IN4(n10), .IN5(
        product[27]), .IN6(n2), .Q(updated_product[2]) );
  AND2X1 U20 ( .IN1(N47), .IN2(n9), .Q(updated_product[24]) );
  AO221X1 U21 ( .IN1(product[49]), .IN2(n10), .IN3(N46), .IN4(n9), .IN5(n11), 
        .Q(updated_product[23]) );
  AO222X1 U22 ( .IN1(N45), .IN2(n9), .IN3(n10), .IN4(product[48]), .IN5(
        product[47]), .IN6(n2), .Q(updated_product[22]) );
  AO222X1 U23 ( .IN1(N44), .IN2(n9), .IN3(product[47]), .IN4(n10), .IN5(
        product[46]), .IN6(n2), .Q(updated_product[21]) );
  AO222X1 U24 ( .IN1(N43), .IN2(n9), .IN3(product[46]), .IN4(n10), .IN5(
        product[45]), .IN6(n11), .Q(updated_product[20]) );
  AO222X1 U25 ( .IN1(N24), .IN2(n9), .IN3(product[27]), .IN4(n10), .IN5(
        product[26]), .IN6(n11), .Q(updated_product[1]) );
  AO222X1 U26 ( .IN1(N42), .IN2(n9), .IN3(product[45]), .IN4(n10), .IN5(
        product[44]), .IN6(n11), .Q(updated_product[19]) );
  AO222X1 U27 ( .IN1(N41), .IN2(n9), .IN3(product[44]), .IN4(n10), .IN5(
        product[43]), .IN6(n11), .Q(updated_product[18]) );
  AO222X1 U28 ( .IN1(N40), .IN2(n9), .IN3(product[43]), .IN4(n10), .IN5(
        product[42]), .IN6(n11), .Q(updated_product[17]) );
  AO222X1 U29 ( .IN1(N39), .IN2(n9), .IN3(product[42]), .IN4(n10), .IN5(
        product[41]), .IN6(n11), .Q(updated_product[16]) );
  AO222X1 U30 ( .IN1(N38), .IN2(n9), .IN3(product[41]), .IN4(n10), .IN5(
        product[40]), .IN6(n11), .Q(updated_product[15]) );
  AO222X1 U31 ( .IN1(N37), .IN2(n9), .IN3(product[40]), .IN4(n10), .IN5(
        product[39]), .IN6(n11), .Q(updated_product[14]) );
  AO222X1 U32 ( .IN1(N36), .IN2(n9), .IN3(product[39]), .IN4(n10), .IN5(
        product[38]), .IN6(n11), .Q(updated_product[13]) );
  AO222X1 U33 ( .IN1(N35), .IN2(n9), .IN3(product[38]), .IN4(n10), .IN5(
        product[37]), .IN6(n11), .Q(updated_product[12]) );
  AO222X1 U34 ( .IN1(N34), .IN2(n9), .IN3(product[37]), .IN4(n10), .IN5(
        product[36]), .IN6(n11), .Q(updated_product[11]) );
  AO222X1 U35 ( .IN1(N33), .IN2(n9), .IN3(product[36]), .IN4(n10), .IN5(n11), 
        .IN6(product[35]), .Q(updated_product[10]) );
  AO222X1 U36 ( .IN1(N23), .IN2(n9), .IN3(product[26]), .IN4(n10), .IN5(n11), 
        .IN6(product[25]), .Q(updated_product[0]) );
  AND2X1 U37 ( .IN1(N21), .IN2(n12), .Q(updated_exponent[8]) );
  AO22X1 U38 ( .IN1(n2), .IN2(new_exponent[7]), .IN3(N20), .IN4(n12), .Q(
        updated_exponent[7]) );
  AO22X1 U39 ( .IN1(n2), .IN2(new_exponent[6]), .IN3(N19), .IN4(n12), .Q(
        updated_exponent[6]) );
  AO22X1 U40 ( .IN1(n2), .IN2(new_exponent[5]), .IN3(N18), .IN4(n12), .Q(
        updated_exponent[5]) );
  AO22X1 U41 ( .IN1(n2), .IN2(new_exponent[4]), .IN3(N17), .IN4(n12), .Q(
        updated_exponent[4]) );
  AO22X1 U42 ( .IN1(n2), .IN2(new_exponent[3]), .IN3(N16), .IN4(n12), .Q(
        updated_exponent[3]) );
  AO22X1 U43 ( .IN1(n2), .IN2(new_exponent[2]), .IN3(N15), .IN4(n12), .Q(
        updated_exponent[2]) );
  AO22X1 U44 ( .IN1(n2), .IN2(new_exponent[1]), .IN3(N14), .IN4(n12), .Q(
        updated_exponent[1]) );
  AO22X1 U45 ( .IN1(n2), .IN2(new_exponent[0]), .IN3(N13), .IN4(n12), .Q(
        updated_exponent[0]) );
  NOR3X0 U46 ( .IN1(N7), .IN2(product[25]), .IN3(n13), .QN(n10) );
  AND3X1 U47 ( .IN1(n14), .IN2(n15), .IN3(product[25]), .Q(n9) );
  NOR2X0 U48 ( .IN1(n14), .IN2(N7), .QN(n11) );
  INVX0 U49 ( .INP(n13), .ZN(n14) );
  NOR2X0 U50 ( .IN1(n16), .IN2(product[49]), .QN(n13) );
  INVX0 U51 ( .INP(product[48]), .ZN(n16) );
  INVX0 U52 ( .INP(n15), .ZN(N7) );
  NOR2X0 U53 ( .IN1(new_exponent[8]), .IN2(n17), .QN(n15) );
  MUX21X1 U54 ( .IN1(n18), .IN2(n19), .S(new_exponent[7]), .Q(n17) );
  AND4X1 U55 ( .IN1(n20), .IN2(new_exponent[6]), .IN3(new_exponent[4]), .IN4(
        new_exponent[5]), .Q(n19) );
  AND4X1 U56 ( .IN1(new_exponent[3]), .IN2(new_exponent[2]), .IN3(
        new_exponent[1]), .IN4(new_exponent[0]), .Q(n20) );
  NOR2X0 U57 ( .IN1(n21), .IN2(n22), .QN(n18) );
  OR4X1 U58 ( .IN1(n23), .IN2(new_exponent[0]), .IN3(new_exponent[1]), .IN4(
        new_exponent[2]), .Q(n22) );
  AND4X1 U59 ( .IN1(n24), .IN2(n25), .IN3(n26), .IN4(n27), .Q(n23) );
  NOR4X0 U60 ( .IN1(n28), .IN2(product[42]), .IN3(product[44]), .IN4(
        product[43]), .QN(n27) );
  OR3X1 U61 ( .IN1(product[46]), .IN2(product[47]), .IN3(product[45]), .Q(n28)
         );
  NOR4X0 U62 ( .IN1(n29), .IN2(product[36]), .IN3(product[38]), .IN4(
        product[37]), .QN(n26) );
  OR3X1 U63 ( .IN1(product[40]), .IN2(product[41]), .IN3(product[39]), .Q(n29)
         );
  NOR4X0 U64 ( .IN1(n30), .IN2(product[30]), .IN3(product[32]), .IN4(
        product[31]), .QN(n25) );
  OR3X1 U65 ( .IN1(product[34]), .IN2(product[35]), .IN3(product[33]), .Q(n30)
         );
  NOR4X0 U66 ( .IN1(n31), .IN2(product[27]), .IN3(product[29]), .IN4(
        product[28]), .QN(n24) );
  OR2X1 U67 ( .IN1(product[25]), .IN2(product[26]), .Q(n31) );
  OR4X1 U68 ( .IN1(new_exponent[3]), .IN2(new_exponent[4]), .IN3(
        new_exponent[5]), .IN4(new_exponent[6]), .Q(n21) );
endmodule


module normalize2_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(SUM[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module normalize2_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[8]), .IN2(A[8]), .Q(SUM[8]) );
endmodule


module normalize2 ( clk, reset, updated_product, updated_exponent, 
        final_product_o, final_exponent_o, exception2_o, new_sign, new_sign2, 
        exception1, exception12, add_r, add_exception_1, add_r2, 
        add_exception_2, s, s2 );
  input [24:0] updated_product;
  input [8:0] updated_exponent;
  output [24:0] final_product_o;
  output [8:0] final_exponent_o;
  input [31:0] add_r;
  output [31:0] add_r2;
  input clk, reset, new_sign, exception1, add_exception_1, s;
  output exception2_o, new_sign2, exception12, add_exception_2, s2;
  wire   N7, N13, N14, N15, N16, N17, N18, N19, N20, N21, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31;
  wire   [8:0] final_exponent;
  wire   [24:0] final_product;

  DFFARX1 add_exception_2_reg ( .D(add_exception_1), .CLK(clk), .RSTB(n8), .Q(
        add_exception_2) );
  DFFARX1 s2_reg ( .D(s), .CLK(clk), .RSTB(n8), .Q(s2) );
  DFFARX1 \final_exponent_o_reg[8]  ( .D(final_exponent[8]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[8]) );
  DFFARX1 \final_exponent_o_reg[7]  ( .D(final_exponent[7]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[7]) );
  DFFARX1 \final_exponent_o_reg[6]  ( .D(final_exponent[6]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[6]) );
  DFFARX1 \final_exponent_o_reg[5]  ( .D(final_exponent[5]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[5]) );
  DFFARX1 \final_exponent_o_reg[4]  ( .D(final_exponent[4]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[4]) );
  DFFARX1 \final_exponent_o_reg[3]  ( .D(final_exponent[3]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[3]) );
  DFFARX1 \final_exponent_o_reg[2]  ( .D(final_exponent[2]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[2]) );
  DFFARX1 \final_exponent_o_reg[1]  ( .D(final_exponent[1]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[1]) );
  DFFARX1 \final_exponent_o_reg[0]  ( .D(final_exponent[0]), .CLK(clk), .RSTB(
        n8), .Q(final_exponent_o[0]) );
  DFFARX1 \final_product_o_reg[24]  ( .D(final_product[24]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[24]) );
  DFFARX1 \final_product_o_reg[23]  ( .D(final_product[23]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[23]) );
  DFFARX1 \final_product_o_reg[22]  ( .D(final_product[22]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[22]) );
  DFFARX1 \final_product_o_reg[21]  ( .D(final_product[21]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[21]) );
  DFFARX1 \final_product_o_reg[20]  ( .D(final_product[20]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[20]) );
  DFFARX1 \final_product_o_reg[19]  ( .D(final_product[19]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[19]) );
  DFFARX1 \final_product_o_reg[18]  ( .D(final_product[18]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[18]) );
  DFFARX1 \final_product_o_reg[17]  ( .D(final_product[17]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[17]) );
  DFFARX1 \final_product_o_reg[16]  ( .D(final_product[16]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[16]) );
  DFFARX1 \final_product_o_reg[15]  ( .D(final_product[15]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[15]) );
  DFFARX1 \final_product_o_reg[14]  ( .D(final_product[14]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[14]) );
  DFFARX1 \final_product_o_reg[13]  ( .D(final_product[13]), .CLK(clk), .RSTB(
        n7), .Q(final_product_o[13]) );
  DFFARX1 \final_product_o_reg[12]  ( .D(final_product[12]), .CLK(clk), .RSTB(
        n6), .Q(final_product_o[12]) );
  DFFARX1 \final_product_o_reg[11]  ( .D(final_product[11]), .CLK(clk), .RSTB(
        n6), .Q(final_product_o[11]) );
  DFFARX1 \final_product_o_reg[10]  ( .D(final_product[10]), .CLK(clk), .RSTB(
        n6), .Q(final_product_o[10]) );
  DFFARX1 \final_product_o_reg[9]  ( .D(final_product[9]), .CLK(clk), .RSTB(n6), .Q(final_product_o[9]) );
  DFFARX1 \final_product_o_reg[8]  ( .D(final_product[8]), .CLK(clk), .RSTB(n6), .Q(final_product_o[8]) );
  DFFARX1 \final_product_o_reg[7]  ( .D(final_product[7]), .CLK(clk), .RSTB(n6), .Q(final_product_o[7]) );
  DFFARX1 \final_product_o_reg[6]  ( .D(final_product[6]), .CLK(clk), .RSTB(n6), .Q(final_product_o[6]) );
  DFFARX1 \final_product_o_reg[5]  ( .D(final_product[5]), .CLK(clk), .RSTB(n6), .Q(final_product_o[5]) );
  DFFARX1 \final_product_o_reg[4]  ( .D(final_product[4]), .CLK(clk), .RSTB(n6), .Q(final_product_o[4]) );
  DFFARX1 \final_product_o_reg[3]  ( .D(final_product[3]), .CLK(clk), .RSTB(n6), .Q(final_product_o[3]) );
  DFFARX1 \final_product_o_reg[2]  ( .D(final_product[2]), .CLK(clk), .RSTB(n6), .Q(final_product_o[2]) );
  DFFARX1 \final_product_o_reg[1]  ( .D(final_product[1]), .CLK(clk), .RSTB(n6), .Q(final_product_o[1]) );
  DFFARX1 \final_product_o_reg[0]  ( .D(final_product[0]), .CLK(clk), .RSTB(n5), .Q(final_product_o[0]) );
  DFFARX1 exception2_o_reg ( .D(N7), .CLK(clk), .RSTB(n5), .Q(exception2_o) );
  DFFARX1 new_sign2_reg ( .D(new_sign), .CLK(clk), .RSTB(n5), .Q(new_sign2) );
  DFFARX1 exception12_reg ( .D(exception1), .CLK(clk), .RSTB(n5), .Q(
        exception12) );
  DFFARX1 \add_r2_reg[31]  ( .D(add_r[31]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[31]) );
  DFFARX1 \add_r2_reg[30]  ( .D(add_r[30]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[30]) );
  DFFARX1 \add_r2_reg[29]  ( .D(add_r[29]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[29]) );
  DFFARX1 \add_r2_reg[28]  ( .D(add_r[28]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[28]) );
  DFFARX1 \add_r2_reg[27]  ( .D(add_r[27]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[27]) );
  DFFARX1 \add_r2_reg[26]  ( .D(add_r[26]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[26]) );
  DFFARX1 \add_r2_reg[25]  ( .D(add_r[25]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[25]) );
  DFFARX1 \add_r2_reg[24]  ( .D(add_r[24]), .CLK(clk), .RSTB(n5), .Q(
        add_r2[24]) );
  DFFARX1 \add_r2_reg[23]  ( .D(add_r[23]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[23]) );
  DFFARX1 \add_r2_reg[22]  ( .D(add_r[22]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[22]) );
  DFFARX1 \add_r2_reg[21]  ( .D(add_r[21]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[21]) );
  DFFARX1 \add_r2_reg[20]  ( .D(add_r[20]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[20]) );
  DFFARX1 \add_r2_reg[19]  ( .D(add_r[19]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[19]) );
  DFFARX1 \add_r2_reg[18]  ( .D(add_r[18]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[18]) );
  DFFARX1 \add_r2_reg[17]  ( .D(add_r[17]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[17]) );
  DFFARX1 \add_r2_reg[16]  ( .D(add_r[16]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[16]) );
  DFFARX1 \add_r2_reg[15]  ( .D(add_r[15]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[15]) );
  DFFARX1 \add_r2_reg[14]  ( .D(add_r[14]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[14]) );
  DFFARX1 \add_r2_reg[13]  ( .D(add_r[13]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[13]) );
  DFFARX1 \add_r2_reg[12]  ( .D(add_r[12]), .CLK(clk), .RSTB(n4), .Q(
        add_r2[12]) );
  DFFARX1 \add_r2_reg[11]  ( .D(add_r[11]), .CLK(clk), .RSTB(n3), .Q(
        add_r2[11]) );
  DFFARX1 \add_r2_reg[10]  ( .D(add_r[10]), .CLK(clk), .RSTB(n3), .Q(
        add_r2[10]) );
  DFFARX1 \add_r2_reg[9]  ( .D(add_r[9]), .CLK(clk), .RSTB(n3), .Q(add_r2[9])
         );
  DFFARX1 \add_r2_reg[8]  ( .D(add_r[8]), .CLK(clk), .RSTB(n3), .Q(add_r2[8])
         );
  DFFARX1 \add_r2_reg[7]  ( .D(add_r[7]), .CLK(clk), .RSTB(n3), .Q(add_r2[7])
         );
  DFFARX1 \add_r2_reg[6]  ( .D(add_r[6]), .CLK(clk), .RSTB(n3), .Q(add_r2[6])
         );
  DFFARX1 \add_r2_reg[5]  ( .D(add_r[5]), .CLK(clk), .RSTB(n3), .Q(add_r2[5])
         );
  DFFARX1 \add_r2_reg[4]  ( .D(add_r[4]), .CLK(clk), .RSTB(n3), .Q(add_r2[4])
         );
  DFFARX1 \add_r2_reg[3]  ( .D(add_r[3]), .CLK(clk), .RSTB(n3), .Q(add_r2[3])
         );
  DFFARX1 \add_r2_reg[2]  ( .D(add_r[2]), .CLK(clk), .RSTB(n3), .Q(add_r2[2])
         );
  DFFARX1 \add_r2_reg[1]  ( .D(add_r[1]), .CLK(clk), .RSTB(n3), .Q(add_r2[1])
         );
  DFFARX1 \add_r2_reg[0]  ( .D(add_r[0]), .CLK(clk), .RSTB(n3), .Q(add_r2[0])
         );
  normalize2_DW01_inc_0 add_92 ( .A({1'b0, updated_product[24:1]}), .SUM({N47, 
        N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        N32, N31, N30, N29, N28, N27, N26, N25, N24, N23}) );
  normalize2_DW01_inc_1 r66 ( .A(updated_exponent), .SUM({N21, N20, N19, N18, 
        N17, N16, N15, N14, N13}) );
  NOR2X0 U3 ( .IN1(n14), .IN2(N7), .QN(n2) );
  OR2X1 U4 ( .IN1(n9), .IN2(n10), .Q(n12) );
  NBUFFX2 U5 ( .INP(reset), .Z(n3) );
  NBUFFX2 U6 ( .INP(reset), .Z(n4) );
  NBUFFX2 U8 ( .INP(reset), .Z(n5) );
  NBUFFX2 U9 ( .INP(reset), .Z(n6) );
  NBUFFX2 U10 ( .INP(reset), .Z(n7) );
  NBUFFX2 U11 ( .INP(reset), .Z(n8) );
  AO222X1 U12 ( .IN1(N32), .IN2(n9), .IN3(updated_product[10]), .IN4(n10), 
        .IN5(updated_product[9]), .IN6(n11), .Q(final_product[9]) );
  AO222X1 U13 ( .IN1(N31), .IN2(n9), .IN3(updated_product[9]), .IN4(n10), 
        .IN5(updated_product[8]), .IN6(n2), .Q(final_product[8]) );
  AO222X1 U14 ( .IN1(N30), .IN2(n9), .IN3(updated_product[8]), .IN4(n10), 
        .IN5(updated_product[7]), .IN6(n2), .Q(final_product[7]) );
  AO222X1 U15 ( .IN1(N29), .IN2(n9), .IN3(updated_product[7]), .IN4(n10), 
        .IN5(updated_product[6]), .IN6(n2), .Q(final_product[6]) );
  AO222X1 U16 ( .IN1(N28), .IN2(n9), .IN3(updated_product[6]), .IN4(n10), 
        .IN5(updated_product[5]), .IN6(n2), .Q(final_product[5]) );
  AO222X1 U17 ( .IN1(N27), .IN2(n9), .IN3(updated_product[5]), .IN4(n10), 
        .IN5(updated_product[4]), .IN6(n2), .Q(final_product[4]) );
  AO222X1 U18 ( .IN1(N26), .IN2(n9), .IN3(updated_product[4]), .IN4(n10), 
        .IN5(updated_product[3]), .IN6(n2), .Q(final_product[3]) );
  AO222X1 U19 ( .IN1(N25), .IN2(n9), .IN3(updated_product[3]), .IN4(n10), 
        .IN5(updated_product[2]), .IN6(n2), .Q(final_product[2]) );
  AND2X1 U20 ( .IN1(N47), .IN2(n9), .Q(final_product[24]) );
  AO221X1 U21 ( .IN1(updated_product[24]), .IN2(n10), .IN3(N46), .IN4(n9), 
        .IN5(n11), .Q(final_product[23]) );
  AO222X1 U22 ( .IN1(N45), .IN2(n9), .IN3(n10), .IN4(updated_product[23]), 
        .IN5(updated_product[22]), .IN6(n2), .Q(final_product[22]) );
  AO222X1 U23 ( .IN1(N44), .IN2(n9), .IN3(updated_product[22]), .IN4(n10), 
        .IN5(updated_product[21]), .IN6(n2), .Q(final_product[21]) );
  AO222X1 U24 ( .IN1(N43), .IN2(n9), .IN3(updated_product[21]), .IN4(n10), 
        .IN5(updated_product[20]), .IN6(n11), .Q(final_product[20]) );
  AO222X1 U25 ( .IN1(N24), .IN2(n9), .IN3(updated_product[2]), .IN4(n10), 
        .IN5(updated_product[1]), .IN6(n11), .Q(final_product[1]) );
  AO222X1 U26 ( .IN1(N42), .IN2(n9), .IN3(updated_product[20]), .IN4(n10), 
        .IN5(updated_product[19]), .IN6(n11), .Q(final_product[19]) );
  AO222X1 U27 ( .IN1(N41), .IN2(n9), .IN3(updated_product[19]), .IN4(n10), 
        .IN5(updated_product[18]), .IN6(n11), .Q(final_product[18]) );
  AO222X1 U28 ( .IN1(N40), .IN2(n9), .IN3(updated_product[18]), .IN4(n10), 
        .IN5(updated_product[17]), .IN6(n11), .Q(final_product[17]) );
  AO222X1 U29 ( .IN1(N39), .IN2(n9), .IN3(updated_product[17]), .IN4(n10), 
        .IN5(updated_product[16]), .IN6(n11), .Q(final_product[16]) );
  AO222X1 U30 ( .IN1(N38), .IN2(n9), .IN3(updated_product[16]), .IN4(n10), 
        .IN5(updated_product[15]), .IN6(n11), .Q(final_product[15]) );
  AO222X1 U31 ( .IN1(N37), .IN2(n9), .IN3(updated_product[15]), .IN4(n10), 
        .IN5(updated_product[14]), .IN6(n11), .Q(final_product[14]) );
  AO222X1 U32 ( .IN1(N36), .IN2(n9), .IN3(updated_product[14]), .IN4(n10), 
        .IN5(updated_product[13]), .IN6(n11), .Q(final_product[13]) );
  AO222X1 U33 ( .IN1(N35), .IN2(n9), .IN3(updated_product[13]), .IN4(n10), 
        .IN5(updated_product[12]), .IN6(n11), .Q(final_product[12]) );
  AO222X1 U34 ( .IN1(N34), .IN2(n9), .IN3(updated_product[12]), .IN4(n10), 
        .IN5(updated_product[11]), .IN6(n11), .Q(final_product[11]) );
  AO222X1 U35 ( .IN1(N33), .IN2(n9), .IN3(updated_product[11]), .IN4(n10), 
        .IN5(n11), .IN6(updated_product[10]), .Q(final_product[10]) );
  AO222X1 U36 ( .IN1(N23), .IN2(n9), .IN3(updated_product[1]), .IN4(n10), 
        .IN5(n11), .IN6(updated_product[0]), .Q(final_product[0]) );
  AND2X1 U37 ( .IN1(N21), .IN2(n12), .Q(final_exponent[8]) );
  AO22X1 U38 ( .IN1(n2), .IN2(updated_exponent[7]), .IN3(N20), .IN4(n12), .Q(
        final_exponent[7]) );
  AO22X1 U39 ( .IN1(n2), .IN2(updated_exponent[6]), .IN3(N19), .IN4(n12), .Q(
        final_exponent[6]) );
  AO22X1 U40 ( .IN1(n2), .IN2(updated_exponent[5]), .IN3(N18), .IN4(n12), .Q(
        final_exponent[5]) );
  AO22X1 U41 ( .IN1(n2), .IN2(updated_exponent[4]), .IN3(N17), .IN4(n12), .Q(
        final_exponent[4]) );
  AO22X1 U42 ( .IN1(n2), .IN2(updated_exponent[3]), .IN3(N16), .IN4(n12), .Q(
        final_exponent[3]) );
  AO22X1 U43 ( .IN1(n2), .IN2(updated_exponent[2]), .IN3(N15), .IN4(n12), .Q(
        final_exponent[2]) );
  AO22X1 U44 ( .IN1(n2), .IN2(updated_exponent[1]), .IN3(N14), .IN4(n12), .Q(
        final_exponent[1]) );
  AO22X1 U45 ( .IN1(n2), .IN2(updated_exponent[0]), .IN3(N13), .IN4(n12), .Q(
        final_exponent[0]) );
  NOR3X0 U46 ( .IN1(N7), .IN2(updated_product[0]), .IN3(n13), .QN(n10) );
  AND3X1 U47 ( .IN1(n14), .IN2(n15), .IN3(updated_product[0]), .Q(n9) );
  NOR2X0 U48 ( .IN1(n14), .IN2(N7), .QN(n11) );
  INVX0 U49 ( .INP(n13), .ZN(n14) );
  NOR2X0 U50 ( .IN1(n16), .IN2(updated_product[24]), .QN(n13) );
  INVX0 U51 ( .INP(updated_product[23]), .ZN(n16) );
  INVX0 U52 ( .INP(n15), .ZN(N7) );
  NOR2X0 U53 ( .IN1(updated_exponent[8]), .IN2(n17), .QN(n15) );
  MUX21X1 U54 ( .IN1(n18), .IN2(n19), .S(updated_exponent[7]), .Q(n17) );
  AND4X1 U55 ( .IN1(n20), .IN2(updated_exponent[6]), .IN3(updated_exponent[4]), 
        .IN4(updated_exponent[5]), .Q(n19) );
  AND4X1 U56 ( .IN1(updated_exponent[3]), .IN2(updated_exponent[2]), .IN3(
        updated_exponent[1]), .IN4(updated_exponent[0]), .Q(n20) );
  NOR2X0 U57 ( .IN1(n21), .IN2(n22), .QN(n18) );
  OR4X1 U58 ( .IN1(n23), .IN2(updated_exponent[0]), .IN3(updated_exponent[1]), 
        .IN4(updated_exponent[2]), .Q(n22) );
  AND4X1 U59 ( .IN1(n24), .IN2(n25), .IN3(n26), .IN4(n27), .Q(n23) );
  NOR4X0 U60 ( .IN1(n28), .IN2(updated_product[4]), .IN3(updated_product[6]), 
        .IN4(updated_product[5]), .QN(n27) );
  OR3X1 U61 ( .IN1(updated_product[8]), .IN2(updated_product[9]), .IN3(
        updated_product[7]), .Q(n28) );
  NOR4X0 U62 ( .IN1(n29), .IN2(updated_product[1]), .IN3(updated_product[21]), 
        .IN4(updated_product[20]), .QN(n26) );
  OR3X1 U63 ( .IN1(updated_product[2]), .IN2(updated_product[3]), .IN3(
        updated_product[22]), .Q(n29) );
  NOR4X0 U64 ( .IN1(n30), .IN2(updated_product[14]), .IN3(updated_product[16]), 
        .IN4(updated_product[15]), .QN(n25) );
  OR3X1 U65 ( .IN1(updated_product[18]), .IN2(updated_product[19]), .IN3(
        updated_product[17]), .Q(n30) );
  NOR4X0 U66 ( .IN1(n31), .IN2(updated_product[11]), .IN3(updated_product[13]), 
        .IN4(updated_product[12]), .QN(n24) );
  OR2X1 U67 ( .IN1(updated_product[0]), .IN2(updated_product[10]), .Q(n31) );
  OR4X1 U68 ( .IN1(updated_exponent[3]), .IN2(updated_exponent[4]), .IN3(
        updated_exponent[5]), .IN4(updated_exponent[6]), .Q(n21) );
endmodule


module result ( clk, reset, final_exponent, final_product, new_sign, r_o, 
        exception1, exception2, exception_o, add_r, add_exception_1, s );
  input [8:0] final_exponent;
  input [24:0] final_product;
  output [31:0] r_o;
  input [31:0] add_r;
  input clk, reset, new_sign, exception1, exception2, add_exception_1, s;
  output exception_o;
  wire   exception, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n1, n2, n24, n25, n26, n27;
  wire   [31:0] r;

  DFFARX1 \r_o_reg[31]  ( .D(r[31]), .CLK(clk), .RSTB(n25), .Q(r_o[31]) );
  DFFARX1 \r_o_reg[30]  ( .D(r[30]), .CLK(clk), .RSTB(n25), .Q(r_o[30]) );
  DFFARX1 \r_o_reg[29]  ( .D(r[29]), .CLK(clk), .RSTB(n25), .Q(r_o[29]) );
  DFFARX1 \r_o_reg[28]  ( .D(r[28]), .CLK(clk), .RSTB(n25), .Q(r_o[28]) );
  DFFARX1 \r_o_reg[27]  ( .D(r[27]), .CLK(clk), .RSTB(n25), .Q(r_o[27]) );
  DFFARX1 \r_o_reg[26]  ( .D(r[26]), .CLK(clk), .RSTB(n25), .Q(r_o[26]) );
  DFFARX1 \r_o_reg[25]  ( .D(r[25]), .CLK(clk), .RSTB(n25), .Q(r_o[25]) );
  DFFARX1 \r_o_reg[24]  ( .D(r[24]), .CLK(clk), .RSTB(n25), .Q(r_o[24]) );
  DFFARX1 \r_o_reg[23]  ( .D(r[23]), .CLK(clk), .RSTB(n25), .Q(r_o[23]) );
  DFFARX1 \r_o_reg[22]  ( .D(r[22]), .CLK(clk), .RSTB(n24), .Q(r_o[22]) );
  DFFARX1 \r_o_reg[21]  ( .D(r[21]), .CLK(clk), .RSTB(n24), .Q(r_o[21]) );
  DFFARX1 \r_o_reg[20]  ( .D(r[20]), .CLK(clk), .RSTB(n24), .Q(r_o[20]) );
  DFFARX1 \r_o_reg[19]  ( .D(r[19]), .CLK(clk), .RSTB(n24), .Q(r_o[19]) );
  DFFARX1 \r_o_reg[18]  ( .D(r[18]), .CLK(clk), .RSTB(n24), .Q(r_o[18]) );
  DFFARX1 \r_o_reg[17]  ( .D(r[17]), .CLK(clk), .RSTB(n24), .Q(r_o[17]) );
  DFFARX1 \r_o_reg[16]  ( .D(r[16]), .CLK(clk), .RSTB(n24), .Q(r_o[16]) );
  DFFARX1 \r_o_reg[15]  ( .D(r[15]), .CLK(clk), .RSTB(n24), .Q(r_o[15]) );
  DFFARX1 \r_o_reg[14]  ( .D(r[14]), .CLK(clk), .RSTB(n24), .Q(r_o[14]) );
  DFFARX1 \r_o_reg[13]  ( .D(r[13]), .CLK(clk), .RSTB(n24), .Q(r_o[13]) );
  DFFARX1 \r_o_reg[12]  ( .D(r[12]), .CLK(clk), .RSTB(n24), .Q(r_o[12]) );
  DFFARX1 \r_o_reg[11]  ( .D(r[11]), .CLK(clk), .RSTB(n24), .Q(r_o[11]) );
  DFFARX1 \r_o_reg[10]  ( .D(r[10]), .CLK(clk), .RSTB(n2), .Q(r_o[10]) );
  DFFARX1 \r_o_reg[9]  ( .D(r[9]), .CLK(clk), .RSTB(n2), .Q(r_o[9]) );
  DFFARX1 \r_o_reg[8]  ( .D(r[8]), .CLK(clk), .RSTB(n2), .Q(r_o[8]) );
  DFFARX1 \r_o_reg[7]  ( .D(r[7]), .CLK(clk), .RSTB(n2), .Q(r_o[7]) );
  DFFARX1 \r_o_reg[6]  ( .D(r[6]), .CLK(clk), .RSTB(n2), .Q(r_o[6]) );
  DFFARX1 \r_o_reg[5]  ( .D(r[5]), .CLK(clk), .RSTB(n2), .Q(r_o[5]) );
  DFFARX1 \r_o_reg[4]  ( .D(r[4]), .CLK(clk), .RSTB(n2), .Q(r_o[4]) );
  DFFARX1 \r_o_reg[3]  ( .D(r[3]), .CLK(clk), .RSTB(n2), .Q(r_o[3]) );
  DFFARX1 \r_o_reg[2]  ( .D(r[2]), .CLK(clk), .RSTB(n2), .Q(r_o[2]) );
  DFFARX1 \r_o_reg[1]  ( .D(r[1]), .CLK(clk), .RSTB(n2), .Q(r_o[1]) );
  DFFARX1 \r_o_reg[0]  ( .D(r[0]), .CLK(clk), .RSTB(n2), .Q(r_o[0]) );
  DFFARX1 exception_o_reg ( .D(exception), .CLK(clk), .RSTB(n2), .Q(
        exception_o) );
  AO22X1 U8 ( .IN1(add_r[9]), .IN2(n26), .IN3(final_product[9]), .IN4(n3), .Q(
        r[9]) );
  AO22X1 U9 ( .IN1(add_r[8]), .IN2(n26), .IN3(final_product[8]), .IN4(n3), .Q(
        r[8]) );
  AO22X1 U10 ( .IN1(add_r[7]), .IN2(n26), .IN3(final_product[7]), .IN4(n3), 
        .Q(r[7]) );
  AO22X1 U11 ( .IN1(add_r[6]), .IN2(n26), .IN3(final_product[6]), .IN4(n3), 
        .Q(r[6]) );
  AO22X1 U12 ( .IN1(add_r[5]), .IN2(n26), .IN3(final_product[5]), .IN4(n3), 
        .Q(r[5]) );
  AO22X1 U13 ( .IN1(add_r[4]), .IN2(n26), .IN3(final_product[4]), .IN4(n3), 
        .Q(r[4]) );
  AO22X1 U14 ( .IN1(add_r[3]), .IN2(n26), .IN3(final_product[3]), .IN4(n3), 
        .Q(r[3]) );
  AO22X1 U15 ( .IN1(add_r[31]), .IN2(n26), .IN3(new_sign), .IN4(n3), .Q(r[31])
         );
  AO22X1 U16 ( .IN1(add_r[30]), .IN2(n26), .IN3(n4), .IN4(final_exponent[7]), 
        .Q(r[30]) );
  AO22X1 U17 ( .IN1(add_r[2]), .IN2(n1), .IN3(final_product[2]), .IN4(n3), .Q(
        r[2]) );
  AO22X1 U18 ( .IN1(add_r[29]), .IN2(n1), .IN3(n4), .IN4(final_exponent[6]), 
        .Q(r[29]) );
  AO22X1 U19 ( .IN1(add_r[28]), .IN2(n26), .IN3(n4), .IN4(final_exponent[5]), 
        .Q(r[28]) );
  AO22X1 U20 ( .IN1(add_r[27]), .IN2(n26), .IN3(n4), .IN4(final_exponent[4]), 
        .Q(r[27]) );
  AO22X1 U21 ( .IN1(add_r[26]), .IN2(n26), .IN3(n4), .IN4(final_exponent[3]), 
        .Q(r[26]) );
  AO22X1 U22 ( .IN1(add_r[25]), .IN2(n26), .IN3(n4), .IN4(final_exponent[2]), 
        .Q(r[25]) );
  AO22X1 U23 ( .IN1(add_r[24]), .IN2(n26), .IN3(n4), .IN4(final_exponent[1]), 
        .Q(r[24]) );
  AO22X1 U24 ( .IN1(add_r[23]), .IN2(n26), .IN3(n4), .IN4(final_exponent[0]), 
        .Q(r[23]) );
  AND2X1 U25 ( .IN1(n5), .IN2(s), .Q(n4) );
  AO22X1 U26 ( .IN1(add_r[22]), .IN2(n26), .IN3(final_product[22]), .IN4(n3), 
        .Q(r[22]) );
  AO22X1 U27 ( .IN1(add_r[21]), .IN2(n26), .IN3(final_product[21]), .IN4(n3), 
        .Q(r[21]) );
  AO22X1 U28 ( .IN1(add_r[20]), .IN2(n26), .IN3(final_product[20]), .IN4(n3), 
        .Q(r[20]) );
  AO22X1 U29 ( .IN1(add_r[1]), .IN2(n26), .IN3(final_product[1]), .IN4(n3), 
        .Q(r[1]) );
  AO22X1 U30 ( .IN1(add_r[19]), .IN2(n1), .IN3(final_product[19]), .IN4(n3), 
        .Q(r[19]) );
  AO22X1 U31 ( .IN1(add_r[18]), .IN2(n1), .IN3(final_product[18]), .IN4(n3), 
        .Q(r[18]) );
  AO22X1 U32 ( .IN1(add_r[17]), .IN2(n1), .IN3(final_product[17]), .IN4(n3), 
        .Q(r[17]) );
  AO22X1 U33 ( .IN1(add_r[16]), .IN2(n1), .IN3(final_product[16]), .IN4(n3), 
        .Q(r[16]) );
  AO22X1 U34 ( .IN1(add_r[15]), .IN2(n1), .IN3(final_product[15]), .IN4(n3), 
        .Q(r[15]) );
  AO22X1 U35 ( .IN1(add_r[14]), .IN2(n1), .IN3(final_product[14]), .IN4(n3), 
        .Q(r[14]) );
  AO22X1 U36 ( .IN1(add_r[13]), .IN2(n1), .IN3(final_product[13]), .IN4(n3), 
        .Q(r[13]) );
  AO22X1 U37 ( .IN1(add_r[12]), .IN2(n1), .IN3(final_product[12]), .IN4(n3), 
        .Q(r[12]) );
  AO22X1 U38 ( .IN1(add_r[11]), .IN2(n1), .IN3(final_product[11]), .IN4(n3), 
        .Q(r[11]) );
  AO22X1 U39 ( .IN1(add_r[10]), .IN2(n1), .IN3(final_product[10]), .IN4(n3), 
        .Q(r[10]) );
  AO22X1 U40 ( .IN1(add_r[0]), .IN2(n1), .IN3(final_product[0]), .IN4(n3), .Q(
        r[0]) );
  NOR4X0 U41 ( .IN1(exception), .IN2(n7), .IN3(final_product[24]), .IN4(
        final_product[23]), .QN(n6) );
  AO22X1 U42 ( .IN1(add_exception_1), .IN2(n1), .IN3(s), .IN4(n8), .Q(
        exception) );
  OR3X1 U43 ( .IN1(exception2), .IN2(exception1), .IN3(n9), .Q(n8) );
  OA22X1 U44 ( .IN1(n11), .IN2(n12), .IN3(n13), .IN4(n14), .Q(n10) );
  NAND4X0 U45 ( .IN1(final_exponent[7]), .IN2(final_exponent[6]), .IN3(
        final_exponent[5]), .IN4(final_exponent[4]), .QN(n14) );
  NAND4X0 U46 ( .IN1(final_exponent[3]), .IN2(final_exponent[2]), .IN3(
        final_exponent[1]), .IN4(final_exponent[0]), .QN(n13) );
  OR4X1 U47 ( .IN1(n27), .IN2(final_exponent[0]), .IN3(final_exponent[1]), 
        .IN4(final_exponent[2]), .Q(n12) );
  NAND4X0 U48 ( .IN1(n15), .IN2(n16), .IN3(n17), .IN4(n18), .QN(n7) );
  NOR4X0 U49 ( .IN1(n19), .IN2(final_product[4]), .IN3(final_product[6]), 
        .IN4(final_product[5]), .QN(n18) );
  OR3X1 U50 ( .IN1(final_product[8]), .IN2(final_product[9]), .IN3(
        final_product[7]), .Q(n19) );
  NOR4X0 U51 ( .IN1(n20), .IN2(final_product[1]), .IN3(final_product[21]), 
        .IN4(final_product[20]), .QN(n17) );
  OR3X1 U52 ( .IN1(final_product[2]), .IN2(final_product[3]), .IN3(
        final_product[22]), .Q(n20) );
  NOR4X0 U53 ( .IN1(n21), .IN2(final_product[14]), .IN3(final_product[16]), 
        .IN4(final_product[15]), .QN(n16) );
  OR3X1 U54 ( .IN1(final_product[18]), .IN2(final_product[19]), .IN3(
        final_product[17]), .Q(n21) );
  NOR4X0 U55 ( .IN1(n22), .IN2(final_product[11]), .IN3(final_product[13]), 
        .IN4(final_product[12]), .QN(n15) );
  OR2X1 U56 ( .IN1(final_product[0]), .IN2(final_product[10]), .Q(n22) );
  OR4X1 U57 ( .IN1(final_exponent[3]), .IN2(final_exponent[4]), .IN3(n23), 
        .IN4(final_exponent[5]), .Q(n11) );
  OR2X1 U58 ( .IN1(final_exponent[7]), .IN2(final_exponent[6]), .Q(n23) );
  NBUFFX2 U3 ( .INP(n26), .Z(n1) );
  NOR2X0 U4 ( .IN1(n6), .IN2(exception), .QN(n5) );
  NBUFFX2 U5 ( .INP(reset), .Z(n2) );
  NBUFFX2 U6 ( .INP(reset), .Z(n24) );
  NBUFFX2 U7 ( .INP(reset), .Z(n25) );
  NOR2X0 U59 ( .IN1(final_exponent[8]), .IN2(n10), .QN(n9) );
  INVX0 U60 ( .INP(s), .ZN(n26) );
  OA21X1 U61 ( .IN1(n6), .IN2(n5), .IN3(s), .Q(n3) );
  INVX0 U62 ( .INP(n7), .ZN(n27) );
endmodule


module topdut ( a, b, s, clk, reset, r, exception );
  input [31:0] a;
  input [31:0] b;
  output [31:0] r;
  input s, clk, reset;
  output exception;
  wire   new_sign, add_zero_flag, add_greater_flag, add_lesser_flag,
         add_sign_a2, add_sign_b2, s2, new_sign2, add_sign_a3, add_sign_b3, s3,
         add_greater_flag2, new_sign3, new_add_sign, add_sign_a4, add_sign_b4,
         s4, new_sign4, add_exception1, add_exception2, new_add_sign2,
         add_sign_a5, add_sign_b5, s5, new_sign5, add_exception3,
         new_add_sign3, add_exception12, add_exception22, s6, new_sign6,
         add_exception_1, s7, new_sign7, add_exception_2, s8, new_sign8,
         add_exception_3, s9, new_sign9, add_exception_4, s10, new_sign10,
         add_exception_5, s11, new_sign11, add_exception_6, s12, new_sign12,
         add_exception_7, s13, new_sign13, add_exception_8, s14, new_sign14,
         add_exception_9, s15, new_sign15, add_exception_10, s16, new_sign16,
         add_exception_11, s17, new_sign17, add_exception_12, s18, new_sign18,
         add_exception_13, s19, new_sign19, add_exception_14, s20, new_sign20,
         add_exception_15, s21, new_sign21, add_exception_16, s22, new_sign22,
         add_exception_17, s23, new_sign23, add_exception_18, s24, new_sign24,
         add_exception_19, s25, new_sign25, add_exception_20, s26, new_sign26,
         add_exception_21, s27, exception1, new_sign28, add_exception_22, s28,
         exception2, new_sign29, exception12, add_exception_23, s29, n1, n2,
         n3, n4, net50730, net50731, net50732, net50733;
  wire   [8:0] new_exponent;
  wire   [24:0] combined_a;
  wire   [24:0] combined_b;
  wire   [24:0] combined_negative_b;
  wire   [7:0] add_difference;
  wire   [22:0] add_fraction_a2;
  wire   [22:0] add_fraction_b2;
  wire   [7:0] add_exponent_a2;
  wire   [50:0] product1;
  wire   [24:0] combined_b2;
  wire   [24:0] combined_negative_b2;
  wire   [8:0] new_exponent2;
  wire   [23:0] add_combined_a;
  wire   [23:0] add_combined_b;
  wire   [7:0] new_add_exponent;
  wire   [50:0] product2;
  wire   [24:0] combined_b3;
  wire   [24:0] combined_negative_b3;
  wire   [8:0] new_exponent3;
  wire   [24:0] add_sum;
  wire   [7:0] new_add_exponent2;
  wire   [50:0] product3;
  wire   [24:0] combined_b4;
  wire   [24:0] combined_negative_b4;
  wire   [8:0] new_exponent4;
  wire   [7:0] updated_add_exponent;
  wire   [24:0] updated_add_sum;
  wire   [50:0] product4;
  wire   [24:0] combined_b5;
  wire   [24:0] combined_negative_b5;
  wire   [8:0] new_exponent5;
  wire   [7:0] final_add_exponent;
  wire   [24:0] final_add_sum;
  wire   [50:0] product5;
  wire   [24:0] combined_b6;
  wire   [24:0] combined_negative_b6;
  wire   [8:0] new_exponent6;
  wire   [31:0] add_r;
  wire   [50:0] product6;
  wire   [24:0] combined_b7;
  wire   [24:0] combined_negative_b7;
  wire   [8:0] new_exponent7;
  wire   [31:0] add_r2;
  wire   [50:0] product7;
  wire   [24:0] combined_b8;
  wire   [24:0] combined_negative_b8;
  wire   [8:0] new_exponent8;
  wire   [31:0] add_r3;
  wire   [50:0] product8;
  wire   [24:0] combined_b9;
  wire   [24:0] combined_negative_b9;
  wire   [8:0] new_exponent9;
  wire   [31:0] add_r4;
  wire   [50:0] product9;
  wire   [24:0] combined_b10;
  wire   [24:0] combined_negative_b10;
  wire   [8:0] new_exponent10;
  wire   [31:0] add_r5;
  wire   [50:0] product10;
  wire   [24:0] combined_b11;
  wire   [24:0] combined_negative_b11;
  wire   [8:0] new_exponent11;
  wire   [31:0] add_r6;
  wire   [50:0] product11;
  wire   [24:0] combined_b12;
  wire   [24:0] combined_negative_b12;
  wire   [8:0] new_exponent12;
  wire   [31:0] add_r7;
  wire   [50:0] product12;
  wire   [24:0] combined_b13;
  wire   [24:0] combined_negative_b13;
  wire   [8:0] new_exponent13;
  wire   [31:0] add_r8;
  wire   [50:0] product13;
  wire   [24:0] combined_b14;
  wire   [24:0] combined_negative_b14;
  wire   [8:0] new_exponent14;
  wire   [31:0] add_r9;
  wire   [50:0] product14;
  wire   [24:0] combined_b15;
  wire   [24:0] combined_negative_b15;
  wire   [8:0] new_exponent15;
  wire   [31:0] add_r10;
  wire   [50:0] product15;
  wire   [24:0] combined_b16;
  wire   [24:0] combined_negative_b16;
  wire   [8:0] new_exponent16;
  wire   [31:0] add_r11;
  wire   [50:0] product16;
  wire   [24:0] combined_b17;
  wire   [24:0] combined_negative_b17;
  wire   [8:0] new_exponent17;
  wire   [31:0] add_r12;
  wire   [50:0] product17;
  wire   [24:0] combined_b18;
  wire   [24:0] combined_negative_b18;
  wire   [8:0] new_exponent18;
  wire   [31:0] add_r13;
  wire   [50:0] product18;
  wire   [24:0] combined_b19;
  wire   [24:0] combined_negative_b19;
  wire   [8:0] new_exponent19;
  wire   [31:0] add_r14;
  wire   [50:0] product19;
  wire   [24:0] combined_b20;
  wire   [24:0] combined_negative_b20;
  wire   [8:0] new_exponent20;
  wire   [31:0] add_r15;
  wire   [50:0] product20;
  wire   [24:0] combined_b21;
  wire   [24:0] combined_negative_b21;
  wire   [8:0] new_exponent21;
  wire   [31:0] add_r16;
  wire   [50:0] product21;
  wire   [24:0] combined_b22;
  wire   [24:0] combined_negative_b22;
  wire   [8:0] new_exponent22;
  wire   [31:0] add_r17;
  wire   [50:0] product22;
  wire   [24:0] combined_b23;
  wire   [24:0] combined_negative_b23;
  wire   [8:0] new_exponent23;
  wire   [31:0] add_r18;
  wire   [50:0] product23;
  wire   [24:0] combined_b24;
  wire   [24:0] combined_negative_b24;
  wire   [8:0] new_exponent24;
  wire   [31:0] add_r19;
  wire   [50:0] product24;
  wire   [24:0] combined_b25;
  wire   [24:0] combined_negative_b25;
  wire   [8:0] new_exponent25;
  wire   [31:0] add_r20;
  wire   [50:0] product25;
  wire   [8:0] new_exponent26;
  wire   [31:0] add_r21;
  wire   [8:0] updated_exponent;
  wire   [24:0] updated_product;
  wire   [31:0] add_r22;
  wire   [24:0] final_product;
  wire   [8:0] final_exponent;
  wire   [31:0] add_r23;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53;

  combined c1 ( .clk(clk), .reset(n1), .exponent_a(a[30:23]), .exponent_b(
        b[30:23]), .fraction_a(a[22:0]), .fraction_b(b[22:0]), .sign_a(a[31]), 
        .sign_b(b[31]), .new_sign_o(new_sign), .new_exponent_o(new_exponent), 
        .combined_a_o({SYNOPSYS_UNCONNECTED__0, combined_a[23:0]}), 
        .combined_b_o({SYNOPSYS_UNCONNECTED__1, combined_b[23:0]}), 
        .combined_negative_b_o(combined_negative_b), .add_exponent_a(a[30:23]), 
        .add_exponent_b(b[30:23]), .add_difference_o(add_difference), 
        .add_zero_flag_o(add_zero_flag), .add_greater_flag_o(add_greater_flag), 
        .add_lesser_flag_o(add_lesser_flag), .add_sign_a(a[31]), .add_sign_b(
        b[31]), .add_sign_a2(add_sign_a2), .add_sign_b2(add_sign_b2), 
        .add_fraction_a(a[22:0]), .add_fraction_b(b[22:0]), .add_fraction_a2(
        add_fraction_a2), .add_fraction_b2(add_fraction_b2), .add_exponent_a2(
        add_exponent_a2), .s(s), .s2(s2) );
  booth b1 ( .clk(clk), .reset(n4), .combined_a({net50732, combined_a[23:0]}), 
        .combined_b({net50733, combined_b[23:0]}), .combined_negative_b(
        combined_negative_b), .product_o({product1[50:1], 
        SYNOPSYS_UNCONNECTED__2}), .combined_b2({SYNOPSYS_UNCONNECTED__3, 
        combined_b2[23:0]}), .combined_negative_b2(combined_negative_b2), 
        .new_exponent(new_exponent), .new_exponent2(new_exponent2), .new_sign(
        new_sign), .new_sign2(new_sign2), .add_exponent_a(add_exponent_a2), 
        .add_difference(add_difference), .add_zero_flag(add_zero_flag), 
        .add_greater_flag(add_greater_flag), .add_lesser_flag(add_lesser_flag), 
        .add_fraction_a(add_fraction_a2), .add_fraction_b(add_fraction_b2), 
        .add_combined_a_o(add_combined_a), .add_combined_b_o(add_combined_b), 
        .new_add_exponent_o(new_add_exponent), .add_sign_a2(add_sign_a2), 
        .add_sign_b2(add_sign_b2), .add_sign_a3(add_sign_a3), .add_sign_b3(
        add_sign_b3), .s(s2), .s2(s3), .add_greater_flag2(add_greater_flag2)
         );
  booth2 b2 ( .clk(clk), .reset(n1), .product1({product1[50:1], 1'b0}), 
        .combined_b({net50731, combined_b2[23:0]}), .combined_negative_b(
        combined_negative_b2), .product2_o({product2[50:1], 
        SYNOPSYS_UNCONNECTED__4}), .combined_b2(combined_b3), 
        .combined_negative_b2(combined_negative_b3), .new_exponent(
        new_exponent2), .new_exponent2(new_exponent3), .new_sign(new_sign2), 
        .new_sign2(new_sign3), .add_sign_a(add_sign_a3), .add_sign_b(
        add_sign_b3), .add_new_a(add_combined_a), .add_new_b(add_combined_b), 
        .add_sum_o(add_sum), .add_new_add_sign_o(new_add_sign), .add_sign_a3(
        add_sign_a4), .add_sign_b3(add_sign_b4), .add_new_exponent(
        new_add_exponent), .add_new_exponent2(new_add_exponent2), .s(s3), .s2(
        s4), .add_greater_flag2(add_greater_flag2) );
  booth3 b3 ( .clk(clk), .reset(n1), .product1({product2[50:1], 1'b0}), 
        .combined_b(combined_b3), .combined_negative_b(combined_negative_b3), 
        .product2_o({product3[50:1], SYNOPSYS_UNCONNECTED__5}), .combined_b2(
        combined_b4), .combined_negative_b2(combined_negative_b4), 
        .new_exponent(new_exponent3), .new_exponent2(new_exponent4), 
        .new_sign(new_sign3), .new_sign2(new_sign4), .add_sign_a(add_sign_a4), 
        .add_sign_b(add_sign_b4), .add_sum(add_sum), .add_new_exponent(
        new_add_exponent2), .add_updated_exponent_o(updated_add_exponent), 
        .add_updated_add_sum_o(updated_add_sum), .add_exception1_o(
        add_exception1), .add_exception2_o(add_exception2), .add_new_sign(
        new_add_sign), .add_new_sign2(new_add_sign2), .add_sign_a5(add_sign_a5), .add_sign_b5(add_sign_b5), .s(s4), .s2(s5) );
  booth4 b4 ( .clk(clk), .reset(n1), .product1({product3[50:1], 1'b0}), 
        .combined_b(combined_b4), .combined_negative_b(combined_negative_b4), 
        .product2_o({product4[50:1], SYNOPSYS_UNCONNECTED__6}), .combined_b2(
        combined_b5), .combined_negative_b2(combined_negative_b5), 
        .new_exponent(new_exponent4), .new_exponent2(new_exponent5), 
        .new_sign(new_sign4), .new_sign2(new_sign5), .add_sign_a(add_sign_a5), 
        .add_sign_b(add_sign_b5), .add_updated_sum(updated_add_sum), 
        .add_updated_exponent(updated_add_exponent), .add_final_exponent_o(
        final_add_exponent), .add_final_sum_o(final_add_sum), 
        .add_exception3_o(add_exception3), .add_new_sign2(new_add_sign2), 
        .add_new_sign3(new_add_sign3), .add_exception1(add_exception1), 
        .add_exception2(add_exception2), .add_exception12(add_exception12), 
        .add_exception22(add_exception22), .s(s5), .s2(s6) );
  booth5 b5 ( .clk(clk), .reset(reset), .product1({product4[50:1], 1'b0}), 
        .combined_b(combined_b5), .combined_negative_b(combined_negative_b5), 
        .product2_o({product5[50:1], SYNOPSYS_UNCONNECTED__7}), .combined_b2(
        combined_b6), .combined_negative_b2(combined_negative_b6), 
        .new_exponent(new_exponent5), .new_exponent2(new_exponent6), 
        .new_sign(new_sign5), .new_sign2(new_sign6), .add_final_exponent(
        final_add_exponent), .add_final_sum(final_add_sum), .add_new_sign(
        new_add_sign3), .add_r_o(add_r), .add_exception1(add_exception12), 
        .add_exception2(add_exception22), .add_exception3(add_exception3), 
        .add_exception_o(add_exception_1), .s(s6), .s2(s7) );
  booth6_0 b6 ( .clk(clk), .reset(reset), .product1({product5[50:1], 1'b0}), 
        .combined_b(combined_b6), .combined_negative_b(combined_negative_b6), 
        .product2_o({product6[50:1], SYNOPSYS_UNCONNECTED__8}), .combined_b2(
        combined_b7), .combined_negative_b2(combined_negative_b7), 
        .new_exponent(new_exponent6), .new_exponent2(new_exponent7), 
        .new_sign(new_sign6), .new_sign2(new_sign7), .add_r(add_r), 
        .add_exception_1(add_exception_1), .add_r2(add_r2), .add_exception_2(
        add_exception_2), .s(s7), .s2(s8) );
  booth6_19 b7 ( .clk(clk), .reset(n4), .product1({product6[50:1], 1'b0}), 
        .combined_b(combined_b7), .combined_negative_b(combined_negative_b7), 
        .product2_o({product7[50:1], SYNOPSYS_UNCONNECTED__9}), .combined_b2(
        combined_b8), .combined_negative_b2(combined_negative_b8), 
        .new_exponent(new_exponent7), .new_exponent2(new_exponent8), 
        .new_sign(new_sign7), .new_sign2(new_sign8), .add_r(add_r2), 
        .add_exception_1(add_exception_2), .add_r2(add_r3), .add_exception_2(
        add_exception_3), .s(s8), .s2(s9) );
  booth6_18 b8 ( .clk(clk), .reset(n1), .product1({product7[50:1], 1'b0}), 
        .combined_b(combined_b8), .combined_negative_b(combined_negative_b8), 
        .product2_o({product8[50:1], SYNOPSYS_UNCONNECTED__10}), .combined_b2(
        combined_b9), .combined_negative_b2(combined_negative_b9), 
        .new_exponent(new_exponent8), .new_exponent2(new_exponent9), 
        .new_sign(new_sign8), .new_sign2(new_sign9), .add_r(add_r3), 
        .add_exception_1(add_exception_3), .add_r2(add_r4), .add_exception_2(
        add_exception_4), .s(s9), .s2(s10) );
  booth6_17 b9 ( .clk(clk), .reset(n2), .product1({product8[50:1], 1'b0}), 
        .combined_b(combined_b9), .combined_negative_b(combined_negative_b9), 
        .product2_o({product9[50:1], SYNOPSYS_UNCONNECTED__11}), .combined_b2(
        combined_b10), .combined_negative_b2(combined_negative_b10), 
        .new_exponent(new_exponent9), .new_exponent2(new_exponent10), 
        .new_sign(new_sign9), .new_sign2(new_sign10), .add_r(add_r4), 
        .add_exception_1(add_exception_4), .add_r2(add_r5), .add_exception_2(
        add_exception_5), .s(s10), .s2(s11) );
  booth6_16 b10 ( .clk(clk), .reset(n2), .product1({product9[50:1], 1'b0}), 
        .combined_b(combined_b10), .combined_negative_b(combined_negative_b10), 
        .product2_o({product10[50:1], SYNOPSYS_UNCONNECTED__12}), 
        .combined_b2(combined_b11), .combined_negative_b2(
        combined_negative_b11), .new_exponent(new_exponent10), .new_exponent2(
        new_exponent11), .new_sign(new_sign10), .new_sign2(new_sign11), 
        .add_r(add_r5), .add_exception_1(add_exception_5), .add_r2(add_r6), 
        .add_exception_2(add_exception_6), .s(s11), .s2(s12) );
  booth6_15 b11 ( .clk(clk), .reset(n2), .product1({product10[50:1], 1'b0}), 
        .combined_b(combined_b11), .combined_negative_b(combined_negative_b11), 
        .product2_o({product11[50:1], SYNOPSYS_UNCONNECTED__13}), 
        .combined_b2(combined_b12), .combined_negative_b2(
        combined_negative_b12), .new_exponent(new_exponent11), .new_exponent2(
        new_exponent12), .new_sign(new_sign11), .new_sign2(new_sign12), 
        .add_r(add_r6), .add_exception_1(add_exception_6), .add_r2(add_r7), 
        .add_exception_2(add_exception_7), .s(s12), .s2(s13) );
  booth6_14 b12 ( .clk(clk), .reset(n2), .product1({product11[50:1], 1'b0}), 
        .combined_b(combined_b12), .combined_negative_b(combined_negative_b12), 
        .product2_o({product12[50:1], SYNOPSYS_UNCONNECTED__14}), 
        .combined_b2(combined_b13), .combined_negative_b2(
        combined_negative_b13), .new_exponent(new_exponent12), .new_exponent2(
        new_exponent13), .new_sign(new_sign12), .new_sign2(new_sign13), 
        .add_r(add_r7), .add_exception_1(add_exception_7), .add_r2(add_r8), 
        .add_exception_2(add_exception_8), .s(s13), .s2(s14) );
  booth6_13 b13 ( .clk(clk), .reset(n2), .product1({product12[50:1], 1'b0}), 
        .combined_b(combined_b13), .combined_negative_b(combined_negative_b13), 
        .product2_o({product13[50:1], SYNOPSYS_UNCONNECTED__15}), 
        .combined_b2(combined_b14), .combined_negative_b2(
        combined_negative_b14), .new_exponent(new_exponent13), .new_exponent2(
        new_exponent14), .new_sign(new_sign13), .new_sign2(new_sign14), 
        .add_r(add_r8), .add_exception_1(add_exception_8), .add_r2(add_r9), 
        .add_exception_2(add_exception_9), .s(s14), .s2(s15) );
  booth6_12 b14 ( .clk(clk), .reset(n3), .product1({product13[50:1], 1'b0}), 
        .combined_b(combined_b14), .combined_negative_b(combined_negative_b14), 
        .product2_o({product14[50:1], SYNOPSYS_UNCONNECTED__16}), 
        .combined_b2(combined_b15), .combined_negative_b2(
        combined_negative_b15), .new_exponent(new_exponent14), .new_exponent2(
        new_exponent15), .new_sign(new_sign14), .new_sign2(new_sign15), 
        .add_r(add_r9), .add_exception_1(add_exception_9), .add_r2(add_r10), 
        .add_exception_2(add_exception_10), .s(s15), .s2(s16) );
  booth6_11 b15 ( .clk(clk), .reset(n3), .product1({product14[50:1], 1'b0}), 
        .combined_b(combined_b15), .combined_negative_b(combined_negative_b15), 
        .product2_o({product15[50:1], SYNOPSYS_UNCONNECTED__17}), 
        .combined_b2(combined_b16), .combined_negative_b2(
        combined_negative_b16), .new_exponent(new_exponent15), .new_exponent2(
        new_exponent16), .new_sign(new_sign15), .new_sign2(new_sign16), 
        .add_r(add_r10), .add_exception_1(add_exception_10), .add_r2(add_r11), 
        .add_exception_2(add_exception_11), .s(s16), .s2(s17) );
  booth6_10 b16 ( .clk(clk), .reset(n3), .product1({product15[50:1], 1'b0}), 
        .combined_b(combined_b16), .combined_negative_b(combined_negative_b16), 
        .product2_o({product16[50:1], SYNOPSYS_UNCONNECTED__18}), 
        .combined_b2(combined_b17), .combined_negative_b2(
        combined_negative_b17), .new_exponent(new_exponent16), .new_exponent2(
        new_exponent17), .new_sign(new_sign16), .new_sign2(new_sign17), 
        .add_r(add_r11), .add_exception_1(add_exception_11), .add_r2(add_r12), 
        .add_exception_2(add_exception_12), .s(s17), .s2(s18) );
  booth6_9 b17 ( .clk(clk), .reset(n3), .product1({product16[50:1], 1'b0}), 
        .combined_b(combined_b17), .combined_negative_b(combined_negative_b17), 
        .product2_o({product17[50:1], SYNOPSYS_UNCONNECTED__19}), 
        .combined_b2(combined_b18), .combined_negative_b2(
        combined_negative_b18), .new_exponent(new_exponent17), .new_exponent2(
        new_exponent18), .new_sign(new_sign17), .new_sign2(new_sign18), 
        .add_r(add_r12), .add_exception_1(add_exception_12), .add_r2(add_r13), 
        .add_exception_2(add_exception_13), .s(s18), .s2(s19) );
  booth6_8 b18 ( .clk(clk), .reset(n3), .product1({product17[50:1], 1'b0}), 
        .combined_b(combined_b18), .combined_negative_b(combined_negative_b18), 
        .product2_o({product18[50:1], SYNOPSYS_UNCONNECTED__20}), 
        .combined_b2(combined_b19), .combined_negative_b2(
        combined_negative_b19), .new_exponent(new_exponent18), .new_exponent2(
        new_exponent19), .new_sign(new_sign18), .new_sign2(new_sign19), 
        .add_r(add_r13), .add_exception_1(add_exception_13), .add_r2(add_r14), 
        .add_exception_2(add_exception_14), .s(s19), .s2(s20) );
  booth6_7 b19 ( .clk(clk), .reset(n4), .product1({product18[50:1], 1'b0}), 
        .combined_b(combined_b19), .combined_negative_b(combined_negative_b19), 
        .product2_o({product19[50:1], SYNOPSYS_UNCONNECTED__21}), 
        .combined_b2(combined_b20), .combined_negative_b2(
        combined_negative_b20), .new_exponent(new_exponent19), .new_exponent2(
        new_exponent20), .new_sign(new_sign19), .new_sign2(new_sign20), 
        .add_r(add_r14), .add_exception_1(add_exception_14), .add_r2(add_r15), 
        .add_exception_2(add_exception_15), .s(s20), .s2(s21) );
  booth6_6 b20 ( .clk(clk), .reset(n4), .product1({product19[50:1], 1'b0}), 
        .combined_b(combined_b20), .combined_negative_b(combined_negative_b20), 
        .product2_o({product20[50:1], SYNOPSYS_UNCONNECTED__22}), 
        .combined_b2(combined_b21), .combined_negative_b2(
        combined_negative_b21), .new_exponent(new_exponent20), .new_exponent2(
        new_exponent21), .new_sign(new_sign20), .new_sign2(new_sign21), 
        .add_r(add_r15), .add_exception_1(add_exception_15), .add_r2(add_r16), 
        .add_exception_2(add_exception_16), .s(s21), .s2(s22) );
  booth6_5 b21 ( .clk(clk), .reset(n4), .product1({product20[50:1], 1'b0}), 
        .combined_b(combined_b21), .combined_negative_b(combined_negative_b21), 
        .product2_o({product21[50:1], SYNOPSYS_UNCONNECTED__23}), 
        .combined_b2(combined_b22), .combined_negative_b2(
        combined_negative_b22), .new_exponent(new_exponent21), .new_exponent2(
        new_exponent22), .new_sign(new_sign21), .new_sign2(new_sign22), 
        .add_r(add_r16), .add_exception_1(add_exception_16), .add_r2(add_r17), 
        .add_exception_2(add_exception_17), .s(s22), .s2(s23) );
  booth6_4 b22 ( .clk(clk), .reset(n4), .product1({product21[50:1], 1'b0}), 
        .combined_b(combined_b22), .combined_negative_b(combined_negative_b22), 
        .product2_o({product22[50:1], SYNOPSYS_UNCONNECTED__24}), 
        .combined_b2(combined_b23), .combined_negative_b2(
        combined_negative_b23), .new_exponent(new_exponent22), .new_exponent2(
        new_exponent23), .new_sign(new_sign22), .new_sign2(new_sign23), 
        .add_r(add_r17), .add_exception_1(add_exception_17), .add_r2(add_r18), 
        .add_exception_2(add_exception_18), .s(s23), .s2(s24) );
  booth6_3 b23 ( .clk(clk), .reset(reset), .product1({product22[50:1], 1'b0}), 
        .combined_b(combined_b23), .combined_negative_b(combined_negative_b23), 
        .product2_o({product23[50:1], SYNOPSYS_UNCONNECTED__25}), 
        .combined_b2(combined_b24), .combined_negative_b2(
        combined_negative_b24), .new_exponent(new_exponent23), .new_exponent2(
        new_exponent24), .new_sign(new_sign23), .new_sign2(new_sign24), 
        .add_r(add_r18), .add_exception_1(add_exception_18), .add_r2(add_r19), 
        .add_exception_2(add_exception_19), .s(s24), .s2(s25) );
  booth6_2 b24 ( .clk(clk), .reset(reset), .product1({product23[50:1], 1'b0}), 
        .combined_b(combined_b24), .combined_negative_b(combined_negative_b24), 
        .product2_o({product24[50:3], SYNOPSYS_UNCONNECTED__26, product24[1], 
        SYNOPSYS_UNCONNECTED__27}), .combined_b2(combined_b25), 
        .combined_negative_b2(combined_negative_b25), .new_exponent(
        new_exponent24), .new_exponent2(new_exponent25), .new_sign(new_sign24), 
        .new_sign2(new_sign25), .add_r(add_r19), .add_exception_1(
        add_exception_19), .add_r2(add_r20), .add_exception_2(add_exception_20), .s(s25), .s2(s26) );
  booth6_1 b25 ( .clk(clk), .reset(n1), .product1({product24[50:3], net50730, 
        product24[1], 1'b0}), .combined_b(combined_b25), .combined_negative_b(
        combined_negative_b25), .product2_o({SYNOPSYS_UNCONNECTED__28, 
        product25[49:25], SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53}), .new_exponent(new_exponent25), 
        .new_exponent2(new_exponent26), .new_sign(new_sign25), .new_sign2(
        new_sign26), .add_r(add_r20), .add_exception_1(add_exception_20), 
        .add_r2(add_r21), .add_exception_2(add_exception_21), .s(s26), .s2(s27) );
  normalize1 n1_inst ( .clk(clk), .reset(n2), .product({1'b0, product25[49:25], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .new_exponent(new_exponent26), .updated_exponent_o(
        updated_exponent), .updated_product_o(updated_product), .exception_o(
        exception1), .new_sign(new_sign26), .new_sign2(new_sign28), .add_r(
        add_r21), .add_exception_1(add_exception_21), .add_r2(add_r22), 
        .add_exception_2(add_exception_22), .s(s27), .s2(s28) );
  normalize2 n2_inst ( .clk(clk), .reset(n3), .updated_product(updated_product), .updated_exponent(updated_exponent), .final_product_o(final_product), 
        .final_exponent_o(final_exponent), .exception2_o(exception2), 
        .new_sign(new_sign28), .new_sign2(new_sign29), .exception1(exception1), 
        .exception12(exception12), .add_r(add_r22), .add_exception_1(
        add_exception_22), .add_r2(add_r23), .add_exception_2(add_exception_23), .s(s28), .s2(s29) );
  result r2 ( .clk(clk), .reset(n4), .final_exponent(final_exponent), 
        .final_product(final_product), .new_sign(new_sign29), .r_o(r), 
        .exception1(exception12), .exception2(exception2), .exception_o(
        exception), .add_r(add_r23), .add_exception_1(add_exception_23), .s(
        s29) );
  NBUFFX2 U1 ( .INP(reset), .Z(n1) );
  NBUFFX2 U2 ( .INP(reset), .Z(n3) );
  NBUFFX2 U3 ( .INP(reset), .Z(n2) );
  NBUFFX2 U4 ( .INP(reset), .Z(n4) );
endmodule

